`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qsLycJnSmsm2xSPJ6+eF8X2CJ4C2QiTFRc7b5oo0loDjssmNAoem0z5+WKWgk2n+hbvyKwoJKDqt
xZzYwtR++A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KkhmYRpdrcRAjuGoaoAKzHLzxojADYR5u8JWVsdfBY07j8buhUzbqVhyS8W647w+r0viHeoIjKjf
g6HMab5esSqXHpRv5kvF4B9YoXDEeHCFrSkg2fGoYVx73Vq9HlvAWTn6QuoqXU7Zs3eTucKAZS8Q
tHzxQda/csnBDDJsFrE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LVAlIKNVxfqaYW6w8bdLy69mYh9xqAOGiqT9mmX3aiMpbBq5qjWo3SDOVOl2TD+9RNYK1vwcUIlA
puhflk0ZwIXuc048Cg6qBp1t88oxQygWhuhgj8G1RxF970UFW+SVuaha0/w+AZVcc+SXKbKbrZpw
/8pquGt1OwnSSumyQzflNmtZywgj/OUrAZRsuwADg4Xx1lHJb4rlFXbanrm4foXmygKM+0Q1jWEJ
cq52fGmTKDddBuPkpwPpRxFnSQOv/4lWVs6RsULuALHdrDSvAIjJIOgU5QWOVH6GTBWPrAKrRIKu
DlfofrvE4zDiXxvbrEgf5U4yQb6Ay1DER4XzKg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JBIHWWKuV/FwNLzDHe7vf7ZxdIH54GBH/dTVukiZQfQz6LGHf2If2p94tQrhayk8+YXiXuYfkMwJ
wtiUNQQMqkiDsifr0FYJtBJx67siMf8pkn7C23SM2BweiMjv3QSIJUfKOSa3f3mMko44hpojSujz
r+JOCOoR34s4QvCR4h8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A3OAKro0P5A6yC/tfBlIxf3pR4JNeDUcHTDsXQYDUCQON/YwW85ksv5RUFPZaLOI3t2jucdviAeg
y1eNOtWwaQZToWup8Gwo4WhO5yb//ZgSIHbDCEm8fREMVCE0YVOV7BpHTKAtBBaKRLNqgqMSzgno
wGETzVyI9TqaG0q/WO9TkftzshaTTfHMRUXWRss3YZYPoq2owi4naIWnEwTu02BFBt4j5vfOZo9k
zqsFTVebGsaQImouUHT0hiwDw5STlrgMDaEyVA+jSGCkUbUEwoPftIuumG+qpCQ4AQDyGyucyW10
BOl++0osqht+y0fBywObkwlxYrL6FepghOGhaw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bi10pD16jMofRnR8op8scjTh5Hrmwjd6a7SP1XSGEk5AWaCdgXJY8OHae4WPMh+spfC9C2TZJz0J
zfszkjOTkexKhNjA9Uj5OT6WMAVoEjJzHiQ79Q0kmnh6im+Sf7huFf7Nr0Z3BHZihQk42zSyTMF0
WWrI+8N1yroWz9gmBK1pP9PDJc5ZIW1uSpY6xgBFmUAmtOCeUOlTa8kdCh2e5aU1gqhk6NTraQE+
v21r0Z06eH0aTf3RuZJutr0EwUSoTWFLXG68E/PbUbDNyFMGFq+3TAixREGX0BN2wSl1xHA7qn4D
lcwjlRmBczEQpr24sNThtFWLqgKMOWR7Y+5hyg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18016)
`protect data_block
+CwdGzs8KZLjhq+NVu6kq5hPWR1lCtLL2mBB39hdPusBC2MmbIWW37SmHPv5/asvxyZxDg+AgU5w
oZ16Adt0nPGPsZZ/EJfg9ki24nsU861eZDvYf+OBI1L3EimmbWnVSq0uA1kor4+u8v0CFoVNC88Q
UeVZcM7pK+TN591nxWHKr93WHbNqsofwdz5ngK7r1aeRlmbJ3t6e4QilK9QxpEGsARzphF1ZFXiV
/xFO+rwvwm9OjNf/tAzc+xOpX88AFNe2zMZMRrWzuElRuMX4r8WVbGq2/Y76So+D0ETevTA+WoAt
BQ2DBJGtmtFHdMIbWj/c++uswfibShu5Jy7MZ+E0xWOz6YgRkk4RIYJIAZUpgcpG/hd1qUvh3HK5
UIxQVdvUp3cZwP+8+OOXnO/IK61KgZLmLRUuxXFqcEvFF1ZQ4ldGtsIZdltfo23bPShLq8adtnxU
FURnQ40T4m+BA+vZXaBYQ/BBlvyvaOY4CFT/XwYW95uuewttM85cqTowQSaRlTaZpdk2FTcH6HfS
jyz3yyIc/8Bc0Tpqb3FSk2/6uUr9wL96mR8hYKUnlCT8/muOnHcdzEOLKSZTE9fiYo13IjV/lxmz
I4MeooCvJMMxA28/9QKjkklQVs6TLIDJgrdtD/xIBWOpddVVSDIWqhSIv3LnpmVKMWFin2V6Az54
3NUqSicOuxkTxW/nQgkF2scCNYg0Ntz5I2jNKkPoYY62G0tdWwZc7DyqbI10Rf7kTPJpMzg/SmSH
HPG2veRSP1lEzSfIpBkCHTynSZ7Qj0Fa921H3O2VtdlR9Iq/Zgopb5V69laa7+iec8olQmg8iBQY
VslCosxFHLRb+yjBnnZ+YOcq7HD1cdUCh4l6sRX5BsnlU1wyJ3PnV2oE9k4R0+iCg7Td/1817nzl
zZvyFgGMtiRebtDjMZ2dtMmdGXMd6AyrWFf+amkIEMYuCVNwEISF1WAAlEq8aTfgM8tfsSH6Oxuq
kYr4GAq6s9Pvj+jLNuaRnoBb87jG1bd/DYgd76pPizkH+HR4a6bsLcyV9JmvgSoQG8ciYt+Dw/3b
0GadFDSuFCp8TMOwXWrteU+sZqYjARv8ZK4kPgUj2hZW4dBOsBnCHqQWwpxyOEV4iinum9VEtrT+
uut/D0yQuG26++upn7ADkcTH9X2JotWidtKHBPMH/ih7UIU3clUtcldAT7BbJI5rMaYRo0OvRIJ+
sRDENSpKdCxRY6fqmzvsaiXvr2n1pz2SWHiqFvyvxgyQQSKTgKuj/oAOsUFB8bU8R9iSka2gTBsD
CxAuz6w1cKD+yOQDb/1Y+D9iTYVL3qTc+z+yfQrTw7/Zo30E0pChefh8KvXpp6/PY6i27+ejmmDK
QzGbKpt9c6Bftzveruh7scKXlSb2fAfE4eS03MRLMgDCsmzG7tTRQCAdxBWCzfZpF+ENMJWC6Hcb
XfmczX/waoVjDuhOuojs0lkiOna3MBDAB6IbnAndBLpL58tC3a5O2MJqGWsLUGxGNDbahR/p1naC
Y2z3LjC6ChuOJqMK0p0paN4EEEJBnWMhY/6aRnaD+lBB7IXcfln1ZiXOpiOlRbSn6pju4hbEwfWz
y0o8uNxJKaA7lBh2M36Zt97IfghS2zoRpzUgsPDsSE+Is8pPl1qnxPMj2Fu4dzp/hIc7KCi9ZxAK
+saBw4OtE2IUXNJzeLsuAeioXFNKBnVWENzzLBQ84vwTCng2z5Xz5l3IaOB/Oz2aRBjnvLNw85VR
nux+XIm+nXfYW2+YPI0iQzQUxNIde2BOkq2X1zTXCpL0A8EG7F2fNglMUBmd6/T6lr8WzJ6Iy45y
MR6zkTxlKb+3Pw/x9Ew+MvXqLwTDaMK+pELDcURDz7jpD0ojf7ElCphPCXHb0CcQqxeRLUGkQ8WB
TqQI/LsTGfKVtVAs84y9wh3i8w07rao5XPXH8rZU0rBi8N/bCrq8YKJv4rkjcU8cQhhmgvL5fFuC
xOBiJjVlt9h9UUiYJz05JheI/uRQe6/PHmkQD/+H9mVyXcOqE5xNit0kaRt5L6MtRv8W90O9qvCv
UPIRlZTJg6FCKd9wxnNVGkqI9hDwcD/+YdCk2pTAJ2uT8zKoqwSJ43B9FMLb9lFO76yvBJbf7PEL
k9zwhbwV5fhY6kDJpu/RQmA+mvfjyGyw+KkG/xHL4zXI/rY4WqN7i3MIQ/7NXlgo6Qphu1mwgD/M
xBj4XZmIZetVsxv1QDMfJgz6I8XOJ5A//tz15xL2fGlupg++LpB+cfQwklmBsq8rcemC6J4YeOT0
VMjW158hwKhCZhMCQ/m1yEXsrUkqZF7ztdPxg46fzP5Hqi02kLfUxlP44UJixjaqjAyOHQtuVnzX
DhtRlXq5tLVHVNCjGtOiKXtKevG2I3IguUwGAKbxL6zgiKAvFPGXn0ntwfNt+V7TSwZz+7Y0xh13
NuxB3LqXBNq6A/yEz1xMW+ZTaOi8HeB1CNTYqLDUMD71A7D3UAqjnRAtHvO+9De1yQKIa2Bc4iFB
pJLIJ26tnL/gz5puivvxlF71vne0cSCzheg4i5+ijuDAz7i0vZ7/o70WfAnIZo2aHjPZhpiwuCoC
JxXwvuILCaBFFSW1uVgZ8WYVHwZlptCEmd0hD8gPbPaOwFtyXrK3LToV23bZ5Y772C3X2omxY5IV
vLBE9CL/UCTTts/ddX7A0s0Pb5l1I+GPvz4jSmpGRI+n+Lu5O4isl4CJcqr1fewN4E8ooNHskeo/
cqvvqyH5ak4wP8/r5aZoNf+ao8HDIRJtNbrijr+pkpuPYE4bSVF+ae4rPfsarkYWwbOq4+ZG1V2v
hNelSPgVijyJeIuTXKMA8Nv4rFZc3yzAdxEt9e20BeF0P3getkJApB3g8PsRfOgap+CQUo36wZ/v
zqbjeTQpoqqSYHbxoToRU+F66OifJZjEvwmXPGgINvIXvtN/YSbgBZoksbtBwPzcIFtBirgxuRu+
lWTuFrGGLB07dfKH4yRHwNJK2ZuX9UOovzGcKSvxEpXAnEdw6CZ0NmYPuNAp/Z2I9keYzPFKkx/D
OaKFarVZ8SVwrMbd8gYN5cxgHAja8c+4bfwhPtDDzsj0VN5O/ge/guw4rZzB+h6W8O7q6+OQdl8W
b0p+GkaJb7QSRv9FEqOuHNSxCTKh5ED9OI7aELWEK7gLNdO36HXaWL8HZ+Zv3vOQHmn2B1aAvwbi
2aQZguud9Wfhy6sWBlHHuSOZ0/zjVjdz4DI+6nz3zIX1ojTatMCOlQsFC5ykr9UUa8evQ9bUBw62
vTvLQVnQPovG3fQC8G572agXx8pPMRy1lOZo8ewa/p1uSMBvh4GE0e0Ek+Jp+Q247Z0GdaMbUaYt
6DrO/p1VBSWmqWMLoYRcOzKJZdsz3c9Rz8EkWxm7Ew4zOh2V9Jh/sFp95z/ewPU6szUaBrkz/ppL
BJbyg7dNgpDi1So0VE+HZJmE9Avn7hZAleLfeesejVGaPCQOWj4eUuOPB9dTkodAhDXbXb2BA2Ql
4U3kccSOCE6p/u3nhgNZUdbTbKX2/4riq6zV5CEvlMQ2M3E5lEhxRyGczagwMXVIf+frKzKbS+4u
5vh3L8aJEf8+ZXRq0NJiE6JY9PYGenJfxo9SbsF17rLWlngmWOj6h0JwQsOFwtZyuXWDlx7wGAdD
0oZ6vo+1uzddOWJDuBxzMb6DFsq+DcCyLqdq8dYHexNP8IgAgFDYEspB2IG5Zyl9uAVd6f9RFVyq
SPGgV77VZAoQal1B6fKjbMqKUCfUk0VA+39ZRJn/z8vBtLKI/zjYcnG4z72+xLnxLnKXuerGDMUM
W0Fn89ysoTSV9u3aXTyDSEkZ3EFSD932TmyC0godq9I7vGXoUWEYzhvP+ML1HJx3KmlYl0bO9MMm
NvycGw8rcbjw77O+4yPcO6jlem8lmYKtAh4lLXsPQsjc8NjcN+/RCsGKZgQCpj+6mlKeRaEOV65o
WspWClmdeSfs7CUhrpHDgJ67hi6VQ7wfWFx2EcZy74jpApdKvH/O+ZLoK/uRdvjY2KSRI8TcMnNH
/81GEO+EOsRUCEfkgh+6rTytBuK4waQLABfuks3Fu8cmA6Q7Ilfzch0tBGFFV9R2vcVQ5MkfVBtk
XXFDvCEkKNTw70ErfXbV8+o4FY84P5Ux6huV5o/zmeCny/XbfyNBjCh+MpkLzRGWFbhj+3Cx9ZlC
6lHVNO4s9y1D1zOUsqqmX0NV5EYWAcjNufKEe5xsBzgIvEzgA1JPOfpasBo3huaUVGFODt4RshLK
wvFTJZneJMaiflJFkmzj6GcZKJUce+ldPkGqWVQyivqM7q7CvZelya4s6is/hwobjGr1+MSu8QBL
wWmvU5u6C+W5aVLJT3K7LJ+SECR/LrGLhx7GuRnEnwDRcSZrQIuE5gqdGjAwzXSp2AvyHnfun21z
sj7IhUAYPbqDVSNp32vjTtOGsQiMmKO0M6O+vPHchGPFE6XntOesutBPepf13LnFORd8fbd+O8CE
awsruI2HO9MuLjGcSQR9ii6BhiBwjiy37usL0G4uVLONWMK23G8WRYzr75zM28p3ueRR47kIrjrd
vGzrbFZbujy4T5GUafpXir11r9pHI5+qe8xMWbARXwdQvvPILfFofDn0vuMxWChZ2fV8GGxphutk
0QRlnpVpXe3AyFSKQoA4ENGAhAF/CMtE5ZW9MstP0o1+ntLlmpe4sCXt8dfOzy3V/WLL7csuHadN
ir0P/ptt5FSpBXBlPV/OKL2bT/9u6B8hiT7KDuLFNSt4I3aezb1GZ+VyahQFM4N8T4NJlQCF8y61
azUZMYy/xvhsFFDbflCQ6YuhqJ468oNUtJQCovjqh8ZauOZnz90afi173FSSwTiQgJBJY2/caqpW
EoIVlDqDw68OgXcI9KzggiKkcS2mFxsvGoDi7MHMzBmh8JCntBY4vFwH02bhmJkdCIlu8WMg94cV
qirxhnADEyHjkROw/wz9d1V0VEgJpVwhSJhkimS24jutQjLx/x92bh3N3nLQwSy3q8rs17nf2DVU
EyvDVRSoOpwymsUWOlJ1j1168dFIB847lMeM1Jb/oQRBKPfTD+m6/rvrttBiWRNSqdlDhVnvfGxb
G5ClYWKykBvlZZzndotwTOYiXPbiNSBKr87ZpJY98J4vJbmjWqt4E6BDINT3LBSmcaRnShTy2cgf
ywHvgfgWaS3CXzfQ4E1nEjGg80g+bTcDYEFkePM0zk6gsVGotoqw2MZzwQ0mqi53MqxrNq0Fq3kS
KPikOe0U4sPa3jBVcldaMLPFaNSqe2h4ydrp3CPUMGtB6cAzaAQ+c4iL5vZIUMLi4poKMVjbTqz3
WIQTliHJZYhNBkpnVfH1awgwEhvJdH5cr4GZPUG1StOwae5uG7MiqUSALloPe999r2DfzpEoA97R
UR8ZpjkeBP5ALvponfku94jQC7Uj7qKmhtk577G4oDXyUS7f/Gimsw2K7MSECDrit1FrO6EGcdMC
jTEk1QAnVxm34ZIZLoU3XHIDXDWOOfU96dAI0QFrlt47deK8CJIRX0JyXQ99n/juxQpHuqJfYt4/
Eyj2oTiuAgFP0jNuAknTG8HG+R9N+ei19txE+JtV5EWOzC+H3AcVqNldtmhmzHMJwtS07ev+wBjh
rsKwYHBXNVvYw7ztEfhM+B2viXxbxHQbvuay41IIZ0Zn9/Vns8klO3webI8OXSS4jpS/YocVitPj
eVOOV9bMXK+MS+odvgyeqvH9xOhPSQBvVLzhBV8Bl4aBv7QqTBaspRvmcpiXkFbvBdGUhoCS+ei7
UMgKzARga5L1sAk9PSYL1auD7mRYKUqaC/1PhFPgQugLGNxwLDlQqE6NJzwbE0kdkxoo//4xKoYI
OQHqJuz+xdoE38kLLzPZZLn4KqPmO/MkdkH2FtiwWM2VS+DCi38TSlUqg6fF7nQM0/bCZvn2Cj2I
MAJBLargGv8PG65RYYdSBoN3D64FeZ0Sp4ATtIB//5oznIVEe0nJ9Wh27FJSADCCSC1Xl3X2+foI
G6sbiMtHHsaFU78vyq2dOP+JlksVRuukahY983kyzsLXLc4EjiCkLAXN5yKk9hfBB2EsbVLqt8KU
KaftEC9QR57v6dwBDThLH5wIjDTIWb7YFNpOp1zCcKekHTQMiQbP0S2HnGo64tHAtpDVl83OguMV
v1CDaeMU+g0m/w4RLe33T0sOFXRtDFibL+bycz7Ns+7GOVo8Bcyu1TTV3zQDPFwCH3den5mt6k9i
VovF+hliEgmfX/W6orfyPN+Jl+6JLcr4m6IOKO3FQAlb1HkpZ9dCW2ZKVPmrL13pVG1KW2HpG0xA
brHYNduDnBuX+nGX4Mmuz0p1a5h8kBFj9ww6juTsjMuQU9MXSKgq478F0id11Pqh4jTRcXeaKk4b
05Bvzc7jf2nJaB+ScqiqmRmfMLUb+aSHf2iqXSSTa3m9okAH9nH8VMY9M9hAH6OCq6IvgUIFEhe9
UUPH+m1y0UHkiaVZsuyHlqzMK6BgONcctE2YbtZ8AOELl08X4cXoBH8Frn3INnxw+OVpko1Iyb7q
FzZXO0A04eWYt2c0Z14yWJbqvRFOHrRyVBrZAYhG63M+XL7b+gBKsbUOrcv7lEQqPdZnv2X54/Sm
J4JLzTyMyHs7RFIRD8x39Z3lhRXmVvguat11PsFFXlPlOhMExZMZBYDNhCMtSRGwZRug3d17rOVi
eglDi++yJVxaTf4YPamDqvvaXEpgyd+0aHlm3xbKkDf4jm3qbCs8HBWllFmhPDxpUsoqPs9LgKIj
KdAkHen5ffIK4dUkNdEdnEgxzsz+OvJ0mDdx1P8mtPKt6ZJG7gLHCwkuh2vpnLSa360Xl5xuKQja
3SRHFICq218s/PkY2LRDiaFmTmqD62c8ro2oQOgeVp5N2lXhMJjLHcYwdJZ8i7XF8HpfYH+NOYB/
C+IO4ldiYPzORo99i27fvrYOzQ+Ar19a1o015YGD7m2CzhLU+O28u36Q6WXxAK2h/H5OQfYrKeLm
pPgg+eAvjKkM2V6nonRpIzdSIA4hzTTd+w2GJJXbBg5T+T4IphKsrr5di5hdKnf2GLynp7iKjqi3
kxSYbq9shRUbf5UhuCElZEOkJBTNsLBPAhR/WoWOMN7rS9+gvH6uq3buskGECiZf1GEug1hdZNIu
+69u1CB6B919F1SLQ/pN6MhP3cWzNTsVS4/BaOT2ux+02Y4CnWFBxro0897mYwM8hHhiG1rq3rVr
xOZLX+xhU/hUooULblCVzBt1WEpjZyBJUHOHb8vap5tht2yve78uYZLShaRaTwZtNS7VtiyF+6Op
7pU3gbeshYCMNGiefQfaRVaJJcjep4eFLPZ3HbOjndg7a9mhM0XCNOfiA7Z7vNCBA2ZzUVMmX/P4
lGLu8eFep1j6WOQ30bJHFQtaLk8o9HlCOJ6y68d39OJN+ITtiF2Qpt7Mysf+kVYSV6oFSBrXlIBl
YvXlreN6u9i/W55xJuQQPelFd91+HMiLtP85CNsAMta/ZQ2lAdmuTuEg89uVEQqQuKPWwzc3Tnd5
eRtOhCNOkWFeiNs6GabI4xqN/Fiuytf2EfwJjGEjaIEogML8nhrDzhNi0QUep8jazEj9+w9L6yMn
bhq2N1ZMiRzxWygO8TrNChxIxR/gZ0iXuq1+tiMJiuMviscJOccYGNB1Fc9u3+T7NISy7dWxf8kf
6GGKOzoSGewmBXzvCKc29oAe1wCIbuiql5Fzp6RQz+Q0MMVUO0tSUdyM6CnZVt51xrXVSgrHlyyl
XtotavxzXehKhT7xuILprJ/GfgsTGy4kjsYvGski0p44GwIGvugAGLhL0zwReQoZz7wFMG+S/nJL
uAkHtnoHy2nWl+6SjP/z5Dvrw+024KWOFRwwVcDkZzMwheUglQP56VAsENFU3/YutKKP7m+6dIrz
lbJ6e3A/WP8O9KVEfLgwOpA/BsTpx9oEItDZU+KMd945DPutCccrbg+wLAlhaaNKE8PO1xQddlSb
u89uwNz95ionPwB78fw9qDbwmEJcDIxzQrMq5gwb93TnXyHaGfb7wNDDGXWtoR1WHjTYGKGiO+3m
WAqExWv01SJ0yx6y3cWCPpF3XzALZIxLEgnllYA+AujUjWAalM30/C2ITN3m8gtVM+IX7oOqryD5
U5G10XEE1/uNI8eS3kwuMvd9FmhXCLS1rgLNPltWcqW8RCboo8z9AgDy13QL4GgWS4lRoAslsV97
cbCC2vY/yOHUA9Sf2hy5SymB+yXPi9lLcxQx3NJfoOGM0yVVYurxjSs/OVXEaEm9/9T8PrXlFk7S
QasVCtWVIOf3c259YRJ7uSGtc50R+91hL0UNYZLyf6a2EmosywjidHz9w6Y8Cg0B8/souiq1E9DO
9y9GSXncSm58pzh448MynO4fqsutJdb9aAHVtQYYZYOU59HxlvgjhotfVguvz8jWWB6+JLevkQXW
WrF0fjw16nMyr8iB0u+rp/dosIIihpXosj3lQDq9AYBQExvQcwfDTQiUb5AjiFOPmSv6fYFls/Zg
ys+YZEOpH2DKmTNsBBU4Z9bvOflBXhFK3fLt5+m7ENbycILKn2bnxoxXb6036orjPT/5z6HQqMyP
BGzjYi/kXZXklgNkIZROEQ6OOPvGtx3dywSHjvDG3v8Tn2Sb1uPGPXifzKUXwoxZuf/VERehmVMI
1++PT8vyLmGY4SfR1wu/x+kfbKc28sEwsD5IhS9FK4vAv3wAiuNgXRRiFq6U7atSXjV1bOnZMvAX
YZ5TKiGhWpu+BkG9sNMSXzr6VamrNa0Xaa2lRiIZ4Xwro/mchCcdeo/uyxsIwxdh1zPKU4XvtHay
UW9E4tF4TXwl1qaOkrnJCokNt3Kui7UkN2vYKoulT4AfOfKf6/G1N5C7R3WAUNEGhR82/XJdisdx
wWbO0CfEHW13aHiu4vAC24KiPJx+Bu3hIHvRo7lUR+Io2RUaxJiKWd85Jhe5ITlhvuRAO4QN09CE
eZQHsgTMy/VZjyzIqC+OKidZL1X12AjmNSna+wm0YSvEvjU+U41xha0eCLr+i7VpnR9BVCPOxgYy
fJULJXTc9mMmSjmxV4VE9oqdRHD9icvACR/w1b/kmNSOsYoFYahSDyLqcTHxq848h4HDEOx/XKpQ
rGNS+M7RIsc8nOZUvqT9F0mbYmH4jsIJqczmArS8Aotk8JOVFMrdh1VDcG9VVCYc68ZJIPZBBQ2/
nmYGQ0qzTkd7CNvQMClSOb7Lewm6WJ5LIy421kf0jVb8hWRdpIaNOlauhtTna+jsF20mh5zp5mpj
/FoMD4Hiz58t32pawPWAptr6B49o3AwD45H9tcq7EtiyhC4XbTrhgCtlS2249xPJm3P5gT93vtPM
UmHKGkwnVnd7Nk/UQJOYC7i/hDR8H9F6b93xyzFDqGAyCHaOQLfVlTu+5Yq9ljFgw9boFdq8Osho
H0kRbm27kcea6Fxj/USe5UZg+bOr0bHFVV/EqFUhHs0qbmLm5t0UGvyEaRmyJ/Pj6DMDziUQF/iY
MKOT/CcLZ60eZRfM4VPQOGqBiNuk1LxWEQ5XuByfT8dXN6078d5cWomisMNgGHsIsJvSntcNxnJX
cVxbm4MU1P6IaSyFxs0aVssueyLR8dQlzUJx/iSPzWMHgadde6E5BkAU5lJWg4emAIWorAzf0vBn
rC4XvTgYlH3Rf6KNT2DZlbrE3TZu7qKV0zahvOCH8FpJBu9VnDqUB02j75ga8o+MMxG+mPKtQxSi
T3qG3vVErE4iCwgyiFul1w4Eu31LfXgZffVqPju4ZSfpgLzwHBLrdRi/81taxjWnykRrGoWSuWuy
r0v5jC/VQq4FZBN3PPALd6mZMyabecJi8AVzGXRxa+/igbgod9HvpNAb+6pZi8qF0uEbRCood0uy
JvZ4/1jorwHHtCjXkUvMp0XF2hWv+rPwX9fu6WLO727cat5qI0pSnARO4G5Hpj4JAarsATSZ8MOo
AP/n40SPLnDC+W+Kg2dasoGBmOe/gukkfBPlL8ts/jegSPAqlkjZ943lNAi2P6PEveE3sDSahxNo
2r+Uya9XQ9IFR08LNcGDRhhsDS2nPcI9Hq1b4qyzUNeQ5mz7It1GCG66NJoJZtIA16/lkIyzz+IH
z3gLZjBaMLkdZWK0eSQQ9Ff7HSYMz098pSkh6vUTNxt3ZCtVjG7294qb3bLMJS82PI93JMYTe1qX
I+MnIQ8au/CT/rIuQV2SNu154f2mx/Gq85ho+SeEP73rimgOevPm4E/7a7HAbm46YaXHFHACavMs
fBy0LLihcgUIt2d3XNQ7WPk7/s7Ez32pCaCuKLKbKBenOb8LGz3jWvyVYQsIYePhQVHbOCfJqgpX
NErlpymSYZVzip3hGXI+83Ks72dy2y5QDkIJFc8oCorkygTc2D2a5Z8PdoV/RlLwoE6pOPBSAWdZ
RJg2u6WPrj/rDO9TxtQ7oabyhjxz0Am6jjk6w2pTZ22eJTri3+h/QG7jLmkPQnvvAPQuSBzrv2AY
NShTk0iatqFJTlbE9fC4TDR7knPNVs4tf8wUHjBpg3KfTGiLcPMGqV2fNpmWCxrsx/5o62rasvPY
B2aUj6upNIB+SnQ3yG6KuAYx2g/uu96eRlaepSRusB3WLprezXobjy/7BAYR9ouLX/filyGaJMwq
oL6MolPXbKyRM8jwq0YVoKiOXJ6I5JI7pIYO74d3P43FUHTsMknTap00VmJj+DleC/sCbA6JgS5p
kyeWtAyGIPra4AB6mrQusgC+m5teAmoa7rW79LUKjjEM9uRVqxSV6mFB8MqygQp+Kfta/0wLlfhS
meB+/j0XzRe7Q49xSVFako9FNz9s0FkU9ozYH69gIVEs0iP75rcqvfWRSPZ9iD3CP+7xaupR3x55
C2iX132Ny5qmNmmBACrJ3tyU0ItsGA38W044KJzj6SFbQgBOLt9j3spuAulqjndvgNANGEgsoaKX
XxRSnBw9++9Dni0soPFDtR6G7s4wJWLltHFiuqpkLp3e+EiwKawFHt+qXvoTCA/rQhLSfJ67Rk/U
DMicVjHOHnBFTms/G0i8SEyoJaUbD6pOCrCP6rzaAG4L0YY7+NqSvd6zAXLj3mGCd+LC/tjzolpm
NMAVP4nTSUc3Q6Dl8mfSIUBZ8YV+Ugzw9Dp5bvZsr/yZ9L8B2Mi9LPbzWHmzqTa4l6FoJcFrFrzh
yHPZ8dzIdmc72kOotHJ54nGt9y2/+UEKtCPa16orgHbm0j5/Dp66kS1PffiekR3uGohdU6TmzSEM
/3B0K1qFuP9+49Gj+MPkvLdwJpJoW+LBafJ2qmNZEQoVDUL9+RZQ8ViCN0hLBkPQ+PaiIKd1H9Wo
Hde1Chexxf3Ezoal7AfBpVb+C9+Gl2KqEnGhxP8pm3sdsciyLbhaA5rp7U8bAFroAA1lBrCXmN2g
3D/T9jB56rUYJBTIdEBD1C1hZJzKFO7sAB9I6ajhWHhs/GweSkSHSbN+0/t3ztYP4GMNuhEHbXSw
5Aia1Z6iO5/sOJ5a/R4RvojjHVJc3bALCQt8UHNBjks6SCqMV/+rIeG8Rw2oViHyUd+ZiS+iGLup
Vx3UWvzJybhrx9I2coL6dY5KDG5k0BnhO9vNL1VjUveFWuknwoD3+Vd2HbwtgM4skNFEDGuuGgnf
M9LqasMvB008NjxUB4Qwz+9Qt8zPssMpBU3QxQVe3rcZYtVJ8f06NR/SudzH0I/rf4um1XrACsw8
C1Ei/wr4d0oVWYudYivWgFLMPR/LU3yW1ssElXlGNHq9HawQsTMvVjoeNhLuaoeJEoSaEZIshC4A
M6pksHQiqZVJ+bBC+QAAEWkpT7mpXcc7H3j3AUHUFGcuh4nEnZEl5iWBDMkQLyhFfq0Z4+7ytCr8
h5yKKBPM0XNvj4p0qNXCxhKgRn8uIyYHJd6336RTNwFblF3X3XYE/i0yu7BbmoaGY4mw0QfpdLPQ
FXIVne9Ch+hf6FJCDdorZsfo0fMP/+89bxz8ryZ0IqhKiarY6anIAVaiFGoKIUvFO2U4nj04wTHB
XgRKakoQNJ+ljLZb3rCnlM309NXgFeIS2Sakaiatc11W8NsmJTMoyuecfvJqBxOrCz4uNKOuDlz7
g7eusMpuhL+yrZoZFvVBDDS5QRrWNF+u1bUNax/F6D+FBaUNfOjnfwzVEiYQXu10rcHnXFgMtFAr
WiumofpbK6+fokX9xJmSfJppVqrwThqnIAlejvo146OzLILBYJOWeY2a47B0IpQaydZRopJlW7QV
sh1nSudEJrGSYUJFLaz3i8ci63tfThS8GQmd3C/WYS+yAiwFjj2x/e/P9lilbY9y0HWp2/5i6+Ep
UJP3eLYZX/Dc6nintEmJVRCC+m8morA5WiYpEP7CAIg9/2768FybCFX0PwB2j0T2YZbxBCMk+/li
xUpGXoDJ3XBGDl1mXya3r1zMNtR6JtWC0asUDqN6pfORiBP86KLYT4+M/pZfxdAqUfNLyLHKQuLf
V3JCmg16jcwnXh3G6rVXTHkrNh3596pm24wvUkDxfFZpYqAZwvTEgf12gm9u527ueFcAWVBVb6aF
1jTZ865p/PwfH2cWdTTDGWjOPFBEkI9m8AnZR6B99F4Ed5whggVlyOWg7CVD+p14frFHyGIhW0Wi
I9SeQPFoJRCOfCcc6kcAULLpZLM3ntD0fCr6RICiHnEMyO2l+vb6eqqDYIovAc/YRqsQmce4ozCH
vty7/GEotCVm77R1C/OhpPUB2DbSfl7w/JDoLIVJdEolGzdkHNIE3TwXpw5PfbKiaWVGSFFvUdPo
uixH3QjFrrZvT1q8EK5dzY9pC8kUOBEiQB6XvB+tbrKp5PEEptYXiRwZV5oEXnIDDv4g2R1/tU9U
Rm7VE1al/OfdXDdCyvmEuE2g7QMlganZUGKJXLzigfha0ioyq40V3v0/QnYrvbFhBDNMFt1BSacP
gvmyphXV6w+8F7wQIjtLpCTzTk3GrENkiGgd2Ke1jehjeWvjf7Hjn1cuhn2yK2qXa8gPJla6OvkX
PGe+WwBncJmfayeexcFLDv1/biAL5qm/MYD994rocFTUD5HCbCofPdOpI0Cn6Ew9cUxVQbbGcCho
bZRM0BgNwPNL0atiK/arIwilRKbL9w+0jxLfMMR+rO2V6DlsUFZJzA8G9Xm1LiW7Qd2KtkNegoLP
lg4dH3Tu/iJEhizgveZFd+9t8A5X8MfGFc6avN9eh/+hnew2AB3aSXRR2n4RdYdY0va9y15j+bDr
qAcgvhv0R8Qr0GKbESPX/a3Dk6TDRFlbu1BtGZ4r+eZJJwDFyPvDrQS+lqbiQlFIgUuthVO7LMrq
9rn1D+87qfGcoHkwMXHS/agWdfDRz22//iNfPzb8bpU6xk89ZcIoRdIHJXz767MP5Fix31Gtkaw5
+Zeimt1RlzWaXvchZ8Wb/YagVHsQxUt3znp2sPzFNsrooP0NM1OR6kMwKZt1MpamjDMx3OTjxoL8
+cJbPqn1T/GfnulGUKmBfDBkuCRAT5h9TTfp0Bj3fonzTai28k+MWlxdAi5q01UH529sdDVEk/A/
2yTjbFYJI/IndwufnY3C7m4RoagLsPAfWu7o9BuZB7TQTrMz3PJ2zKgunubLv6hxwNxrpJ8++8WJ
KosPLqc9R3kzXQPzVheTIXM0MdGBKWUfJuSGFyw/JKcFYcLnlTRaoPed6qXAGunovyLat/HGKFzV
tUfz/EXS4lhMuG4414wNek8p6ciY58Z7twN5bRwfGlW6glbIOleGxOqkv496+EpSL/lw3rMcNE1M
mzbTfltdlxJ2R9yZu2CnLBZp+v+zWhrmKSGJpIlbIYg1AC6Euxl2M3on3y+RVbH74B94NaEDyZBQ
slm2M7VEaI/eSSI9B0e+xxysergFZYxDshTXUUqtfkgPnpEZPB8zj/Twa8LOmWTIiefwEVx20puA
KoaW6T/FUG4vIRzOQRnrltQjwD/ync1ZtPzKZEcNRBbsUqGTNS7/Y0XHTAoybGSa/z7BuvedEfjS
zfJicMCBQVAdApYISeUminiP60LB+7OjizzevTZj3hoJNL9+5c6qzAsng/aTxRw/snM+yfknrHR5
1j/bh67+J8WYI5nYxATtZRzkdMa8r7QkA9IirAT8IgwGpyx61W9UUq404wloYdiSorxZCdcd5Szp
4TfjGj5+bhHO5YUpy0VhdFD68vlINsvTro4rmLO+tSwWxiTmqC4KRmuaxVospsX1nio21ujO0rB0
E8ImONphUYrO4EM3PpAc8vSr4h0DgVilunjjSeMsJi5p8FYwffrtOMIbMZH/SAfZmX6c4nfdzEox
QvvIROTY7j+9T7iVedstBWinDFN5PgjRUB5CkeGFiUAVYbvrBx3IS6+YofO87eD2stW7//CH9Jmc
p+CpGozXl6teBET4z4Qy9/jKHbPDPEmclSTE4jpnJjzo8ueY+tQB8zUkxz0eb6Lltn+X1pgXvmcQ
Eeq3MyY28TikB0NnsD+EHR3Cj7HYIRMRf6qr4IUgui9rlGSRmfG3wVCZZb/iae6yIIU2+fShjHRD
VQyscF6JYAtfBeYTIveITFWcGoFJEVUWspKtPL/g7TQ+uiOwtR6167wkjprmuTNHAOJSXLmXyeEG
bps4Uh5LLNVLczuDRMRXa9HHzgI7BUJzlxHiahfEvHaUmkPFVzPIHCShi+33xhDg4d2AN+diuyRT
XDGbeB60vn4+H/YLs8fOxQ117xnI0t6+8QegSWJ2hGUs31AVUV+qvlfSioRbT3pLyOErXy1YQSfK
dkI9yY/mvNZNCPFmtChCtO1I5rL57azmiFDM7LUKS19LcRHDly1M507lJpVTSCYwh+kJVWAByyNI
OBYXcUXw9FtC1VpLe6BVMgxPRMkG6rpTsJXOldxQY2kXQiJ95UiCKTIqXyyb6l0uwNavh/YaeGhO
Jlk+EV0Jfjsgh9jP7yC+Xr7HTqdjxb2wDfAMAPKQX0rMlYPTgZKzE7KrgisZB+lMmfQAiY2qSWdb
hArCJQQPzXeiavwqzH1NMcyw5VypFdsLm/veIih3waMpUjNGWqn07IIKB4wIBs1UjTLhoc/lrRtH
Uun5Wa/K9rLzQFEdVIuWuelDeK0rq+6A6HLblSRJcQHUCxKK4PNTbZUBgkgXDrfN01ZazV+z1llM
4PPWM4iOHEeKTebDILQyhhcJJPVyunI7FKzOOKqnxnrhCmblDE9qbEUczDaQSvQ7xjBxivNgElq6
LocCtXEFOoCjUnMI4M/wdp8m1nhz/NDEgzza6QL4vQUJc7SdZQ3hsRrqg3oTLxn/LKpgFp09KamY
GJbgF60lk2Sa58jS5ldxnASqFidnKn+eFqqJ43bDzz2TIPsrDgsjiUmwBu+wMivjUNy3WwwACmDS
ivbH6yIA8aX5603xpsjPU+pM7SxMyQKQNqTiJD0DWe1233ChEPDVtakFhuCpFtWe8CQ0iMiVckFS
BPVmATTunBR9FBwFz3jlBRb1LJNiO1Yj68/rCSRgh3JQSi3MPMysH3ZRu/4AOE0NQ7u9mS6TAgpe
0eLm6DsK9kqZKmplIG9zTGkePGmS5rTkteBSTKiN0H3q/EZyg23HOR4hJOENcZov7TbiMT/yDkio
t3ber3PJKphxAvhA0MjoCndU5fxs7yFWyVN3phrz81rOyzvazf59dPAWZ6IJuk0rsGcNDbgXfHIk
dtJ9DZODpTQOtE52IahCwmps9Qy2aBl9+ItYCR9RYMZuzYznBOVrVz57VI7BKJ/REsoj+Kqt1cgV
tvvsqXD39QbuEapdTgILKj9oKVs8eC6q010F+bOVK4d9yRzmIggQ5CfGVcdXYvi5W2NMOSOzPFpC
efOl5Kxb53yRobrvOiR3g3q1ZaEya6Nd7sebZdWMBnEA5bVVNtlCO29rv52HI6VZgN8DmfKN3Tha
LsUnp6jaONbcKUBN39akFGI0+xML9QQzaZAEFkFK7OIR09Km4zzGUnvVjB/NmyO15XiKwh6gyIps
iVnMrN6CDmheJeIL8XJ0mRa5LGinBVPKNLZFZ/nY6LvfjhMJhzEohVA9l2x9LshrV+c4wI8GLGS+
qsw93O4ITXuHMphIGjZwmhZx5v+cBB3gICV2FvHoFsWOJ+84CoEBgAybXOBwWiRIbDhtbCUZDFKD
lWgFgFl6mpnpUYD3sAR9Gl3KbbrOiAkjMmXzy4eZ4L7RK1ZTOdaCRYHYHpeRc7wWz1LwQKM2yrjb
0duOBqUvdpze75AgFKtSwds2TU7she9LGDiQu9xJ/BOpMOijsytDpx4oBQ7vQne7xoS29wYFnHXV
O+KW/mH80RxBZcCdaYJDhPAfVSMqdNbWk/3jkNGz1/kgCZZHVwjJUTuon4W0vGVdc+gxdhB73eOg
EJ/tMHCOIdJoOYC2nXg/QuBwnwfKFlvzK4uq6/8D5BjAGpR++CstMz4EyMgWjaAKiSTLA4zD4dXj
OXgZNEIlizzGN+km0UzHX8NN/QJGESSrL4Px8YNqmJoLkTciolT9s6EHLqTPrqEr6iqS38gd4C7E
Dayglqx6Tl/Y4AbMRZjNTfZqqG+aApm6IoywzukcfWEqQVzPy5oXfMb4aau/Sm+Wg9O9kB2mVBZZ
JUty9IrgZASpH3GiXC6Lu3s+SnqmF+4NQvspVveLcfdHWkLM2rvqBmDnMj/cysZPj4JLZMqFvJQM
HU3Is7ZN/uR4jidKRpmIUrr49hzoB9JpjzmPBVz47kNT5cnCnk/zRqEa14nq/0N7B/r05geK9J6F
WLiqqmBMRzU/YfadGT+ECGmlDBC/Z/jagNMmx7PdeTrx38EiH+m0kLNzqWdR1ES+NcNMCAD+W4JD
Xo0jztBcL88EcbPlbFntkTQ3ltw6anZ0wM3nccI8nTTBIOjW2GHh4f4A3MfLCKMdNIVX8uNkBVyL
0aliCs5JUI5YOfOP/fcORAsLBqLbF1jGToEC9/YDA0SulYEgylSsA6JPPxhHC5bgq0HIHurt96CV
jurySLTKfd90c+zZ4lESccu0m8ELBo5TFyFAq4arSmJgUB70/Jwmgq0/egTcweqrh4SUOXRc2MgV
yjKKE1VsGC7uj8AbpeFhs/k6yEzhGA8+huLWroHLQRVHNvX2q6S2tk5CvXQbzTFgG+ERqjbSUHlM
H3Kzt8biC77Xg9vSJXQcSmk2GsQ2R3w9vYE/7vtC1Fhn54DGDr4NoUkvo+6ZV5tY84WKhvTrFbGe
rP6HHWBR0ydE87eTLUIWHLJALA2S2t/d09beGZCYp5ZUjeinpN6KluzFKKfrRuyfUKzYsqf/i4/2
xCpJDggeMiR7vxLEC8WBuFyrdRu561tafQJ/bawICqmVsVW7eaF4SPJypmbpHHo5R5ehT/ffp7G1
VTJKJ7pyINz5SwWQyW9GGeRBKWYM190z1rvsNP6FYtYXta01qwt5Qf/0R4N6MenUpRVT/eL9vA1p
+lYjWEvDIMKnNts0p6XzQOfcZ/aI9D0fQDZ19VX/IzPRhR0EBrGo/VZbx4Wp/VTl2b2NDTQ2Zz6V
zPiDTTpdPiOTpMGNJJuja7jvDAR4lJGlNaujU9HuwJadygwLvgLikKZ7D5CH/knGkH+2206h9FPC
Kxx1uJ15XHTj0Qlb6aKyN4co/EEIr4efo5z6y3EOLlcfGu/OEHO+Yfv9Xqw7FohbSVVjxQ2pCtE3
RjQ55y3WylqGKdToS6Z3ZpPtK68qhX3n9hRTWU7njEB+Hx3ETeeYK/EgFZoGoQlBoXLnxbMZJzp7
l+RhTfzAFtEG4bxREtnc2Z+pBgiJXBFg0TtuU0/4nH0hP82wBQ+Thg/7REOnS9HY26yzu3oG6L5+
8UBkqvTJ/XNC6raHPQNsjW3zVRh5UsVyI34d8cfBGs7ij7vusQAqlhY0OylVYYh+1mpS09lE6OA6
WvcfEJXIBfFYde33nohnVm4RNPm2W+YKYdrVqc/c/JseMlor06/ot00hZvbiHy3a7/CCYedGQI43
aG50483g9qybPWpYF2jGgC9uq2+hkNRe1nSHDW2+t4P8PGy7+qFWdeQdNEJZxbsMm4Eoadm9XLCH
wpjonOB9h+aikXd4ff1WpS28bTuZ0OXWVdiFg+JFJRem3boLDrjuE/JoouHr11e8Se5gN8RzC56m
hRL06EVgUdebN8L8pqDzoZ7mziJOAyLJHdKBmuwRe+pSknTQRb77gejCJJPAg8pcYsmZ0vn9ND4G
JiqCH0QxaMacnjGDkpo1+IHC5nagiefUxnrx6PMNSNOiBkFcvR9agWzmkUJUFkCJFVtL9KIyIxy7
+SWdlE6/0lm/tFUtOfYE++0Iboo4FEhx6sB1RUCY1nS1PJq24tXuXwPT6zBGEuB8D3fuE3+jX2VD
G2Q5WR+V4fCYw/E0lq55YJ3bUM0ih6OQxxTsncWWRg/Z80zxaRN05ODG4EIn+XNFToOAxYtW0MBM
N/BUoYjL65B1Rl9sm86jsmRNNSmZ7SYnBsi0hfNmh0PfPPmrB5TXHm4oBaEFiyXaHCq+JySw6NPY
LR9LSWTIhhwfbbInSbiB37W3alBaY5b5cd+YRPJ1xxMhixceHTuEHVm8m61lHR3Lo9Z5OSwG/vbQ
pWrjK68hFtPU6LzbYB263wD8Kagj41zmXPvJ2KodVgVeV9IMSvsc2ZMFFXaaFRjwt0nwRWYOxaiE
1D52MnhmUFTM7sJs4yMQ0gvqt1NtuyMw3XUzqmWYyELW9olMqmRe5pUn4PKSEd+87iWpDu7P51RF
P600iz4DcedJH1Uncy2NkjgHiEhOtsVEw1Db8p9PLtChLXsHlpJ34Hm222YyjHnRZO9UWq8ipX8h
MuVX4CeEblo+KQDQxa+zbdZhGwWfxqpV9rCmKGR5jKblM6A1RdZ+thYqM+6YNfss2ZWhciwxImtC
fYvV11GVBTY0ze8jAUxZlIc8g7BFJn4CYM4HohbOPUMUYb5Wyf2nSl91XzJJxb0gCnJ8wHMH1ILH
cIKs/yfD3Kx6SMYYHZTMurQuiYXdqc7MKyC6tUtc0EgHWlsMabG/Wah8FqKvwXQVhGsir6Cmwxx9
BnFTOXOgjQV67JOMpSjtpgEjJ9V34qu/+rOjfgV+N9SqU2AzyKV4MQgelfTHxNovI9aEg/xaNnPZ
wIJ2CxF2Wmiyo4Yg/uDTE3lYu8EFI6ydlP9ar7YIKj5+UIPNjhnTCnOIqvXYs9+Au0IgHJ1GYzux
nkXFKkQei3NkqQYbPQ7HRMoWKj7+5NQ6eE8RF3fEloAAajAImVyPykei72l62O71V4N2sfld6qJm
R3JMLqZJd6xYFLfTn66d9WPJ2TR07kirvNK/fd9ljsS3jlll02dZrNIOX3IbABNwDqiQ8cnq1zle
ILxWgg9LWCy3mMtZbQtWMpU36if1ZNJD1s43Khg+FdzXPPFSiczUDLsz+DQwi7623kYI2Lrc3IcP
kyW3uMw6xz9bRaM72KnNLqXic/7LAXlJuy9a5051xKJI7a2bXT9KoNcqAA7/l/0G1mQ1z9ZOHlH0
qvJV9ahsqsr06r6c8dX/67KZN+SNekUWIzrCzGGVJlgja3HfiLWq6pmfmOVyHvQnw83qQlEHCgfS
/7zn6o5N1lWFL0JtMC/R02+T1t/5Bfkm/uEoVItBCSuCUApFlGhjg2A2wJoN9Rwk8JV3noq22MBl
n0XgGqjy2ALX4zU9kP5x0Ju9xhJ4bSiQUe4N7OKkAvQV7lLpizDDQEtmFrlygwSl7LFWc+PLAoCx
VaQGst38TPgjqaOXgMAFK5Mj/NlQJLiPfK2cxeyzpMNHSjADUuWoMnZExCcPag6qttsp21vOw/QK
hOKAcJCr+U9fupc1SWFQDjFI8cvpkNPsBDvdEQ2i7Ehxz8qWwJDzhRfl7brQYdbIyPmG1u/guSpr
UOVizUGLjHl+SXlkxLJntJluqh0RbDserW8esCMqu8a731JYdD114LnoiNimdgsbryPDzGpsihvj
WVpARFJ58D6hhGDivmVN2QJOlOOeu4bCB1cuPf/PbdPHeKqXWrOvmunG6/v8dg4mX+DeZN65VO6M
uMBIUJtn44Kdq4uc1EgxC78rhQPnBltKWPiKAb4adiTYbv3B7b/IyRYvgw0LuMTCGYEy7Qb7h9tR
/2EB9eWvwJFv1/qJovFiMXrHJpTFd4IHzH4Xn0LNEEeaekcrEyXB85aVk+2ntyyIkFSDDog8Oqva
eCCvytqSnUOv+MjRj3Qfsw4PuVWU/soVq+smzIXBe/N+628sbSg06Bwga/b7GAQA13tX3GzvxhSb
ZeIHKVkUAnMkuFxlN3//JcIdUThuw8I13J7iyL/EcPBt0eY8wRuSu3qqJYfzriq9eIiip+jnErpR
jqtc+xKP1eACtF4Wqy67qftYgpgC+lDf/ub8IkMYtYeyYpg5KQiZIseGGeZpl5enO1EUIaw/zIhp
pSyHV5o/8RV1TLJ72nlOASVUhxNn/SYKVqZhYolwLU23F9avO7ic4sb1s8VkyqsRprkq3JSIJ+7L
oHkSmcUbHHYtVWN7Rio88X41j+QLfjR8+x3VU5E2OL67NdhQGW5I/pPsWjI31Di7eaNLhB/p8p8V
iKkoJkw7mE/HpY8dXlx4PyeNmotDdcpF6LFgmcPKyJ90RCRdQL4NglNyxhjs8hO6R2uM74nKG1cp
FGy7gcbyVCbnX2z/BBmY6V+sHcYWpx9KilVSYsV9WE4fzBC/NrEl3AaUUuWrqiMZMngvv+KssjaP
hgov91NWLv923Ppb94LkeZZ+tMJ22rwIYpPlWTVitpn83u6ggmQXdLxxEPj+IZRK/helUjuSj3Ps
bihoPZjSVVyB52Dy43um/wg+4d4sbN/c0MEXSsbwHcnaaDP+GL77mZCSYb8a2muVSxFbaN6iiZMN
+Ps3V0CipVtOpqVEmB1QU6DbjAZZABQ1XgaKgjtAHGefYSnfwBOFvmuoriDSpGj8VWEOVDKGAH+N
8DW7nFYzNC8GlepVetQXfe3cTl9f42LHbuUPIp6eHpmL44d8AEVydYIbGKtKZamRU3/wu0ebKdPQ
N6BanWxOmwz+Y+8hAa4lL3GhPhJ9BJQn4jX36FSwsf/FW3+3yebtoOAnnq/rSKZIexUHbWA0rQxD
3yhoarfwdsINbAYZ2psfmZgyX4wRXrNHwJdziBlJWC++h6lL1eXHq47h2Ej70E9vg4jJG11L7X9h
PRLM13xBLEYmVljWz+9ZSUdMyWt8OSeiiOleWFX1xtOFVBxk1EGr8zrDqwmfGkuUak9yKh1G7TZB
NxcYtwGhj7EN7eyJxxzkm9vnlGXYDqvVAjymeTZy/jDKvENcw3iEPvU/M/SVm21WS9yACahH1sBr
M9QRHp0NL+mRkEnqfOz4dX/a7wm/Vcsu79/nVszG/ZkOULwJQkwuyoBG9gKWc3h/crWrNrgDeCJd
7IPxWWx80dTL7hrlAlyj6TWiBrsIohIqkjWMtfmO11y84/RkHrG3IIAhr6Z64XPYPevxvLxjynhl
wgW6aSiZ6Lc2AqZU9EX1ZbntV2rjFVySt6LeCm3mBb2/DBgc1rSbnQO4yRR032A7wdG1MQJehkHO
gRtajq8N+0PviOFX+VZYQqVMerDO0cyWC90RTBFDeo66JH+UtG26vxM0r50q7isgVzaY5wNIC8J9
u+5omyqoaD15J+80P+Qa93XyfXONJbDIT1zLb+XQcS+k761BWkbNOPswnp5p8HgAx1B9ylo+m3v0
pnK2TNbtjxR74iTLx3wkxUX/l1S8O6PRIaSm3ijXFOroqtJfcdTR/8OsLetRbMALqcReQQOuOc2R
/jV3SvZgtUKAI5v1YA99UqFoLMNd+KNodgIO1pwft8nbQdefbvgqtHCJkWz2eoKtcUv1dH1rOAyr
K646JRm23LQbIXr3mO+UqxH7UjbukLxcTeU5elfYOCvc/JYGCRJb9FfUvMt55gyzSmdI7T3KzfT0
nffmVnlB4ezmhIa3A/ZAZ0d7v5Xiuw0NiIlmaj9ms8gNNn/l+nddIh9HOzPcCWYD/3J6a+GezFHW
6BZG6bNiA17hVFtFY+99DjhnvmlCcAlpCY23SFVlVa73C+2abxAEFDv2X/GvCMfVcMuR0vQ9TD6c
KYcVM1+aG3mjKRbXhH00ye6/kJuMQoZN9JK5JWSt6T2HF9f/87FsaLuUknlipkOSK+yCcwK5lten
isK+qFgvY/KlQgFcfjgWARWu2u2LiYWwsNR+KntGMuG+RwHEWxSr2f39H7yDukSjJr5+j00RUdMC
MrQDuK+WKPlx2zwSK1X/paB3NNseLa6ZaXBBNsXDq2dksYf2Y4Mrv3xFcXRaEo55LomipVtz1HVw
do+1UWuaXm58bkTEsEBJrP5jayrm/InUcz2MryYAw53x+0o55KaixvOSAxp8U0UQRZaOVOpM4kx+
oRuA/4jsaUUGLoAmGJ29bN2i5wC7y5YAQkhBSP+orZzCV3++3zwwbnlC3BTAHQoNjW7rItsUvCWD
iLXNCyJx5WwmtvujiaKLDM4Ta/IouYGmZUaCI1NlLsA8qW4pU0mOWtGT3BW1HIOI7o7T3NAPhI/A
rqe4ph6oF+aafXNqqJKswoENhbNzkG6nUM4dUccn8ZeEzLT4P+DItwgZrPeCKHGBf/AioO+r0xV9
U8AaHBwsSI6Tk9r7/o5JCINxJ5SSeiKXY35PYhfs3UfyRTtc3Xe8xDrc0h0i7fE/1FtLY+HXobqg
iSkE2Rtm70S9/Q0tPKZpaFFrNseC8tdjA4ABWIPrDa0pNvYVHQ3CH77EraE51BDhVK01J7PFleLN
KWblNo7z9duN4hZ0heWfBad4RgnWqT2XnVN97qVpEqcQ5M5EO/2qJg1QKhxQ1A90ZhoOVF/VDzJS
NdF1ZPl9t6qdofp4JwJpRfrKiDzyjbLocz064V42EZ8grkTZQJ7HUfPiZTs4fAieoasdkqziWEr5
k9zg2TMeUfA6+YO0IOc2pgSpoco79zDGEKv+jgRzZCLJDjyA2NHP3UPCv6S6FvCtgJtq8mom/gw2
ZK+npXuHc8eei19XZ1LjiQ/Z+tkEqJhnkHgxWfSpBHct3fCocRY8haQH6adRvU2pa2/iLB+WasgO
rjCilReW2hEtwUr8Zg4w7AKVsf0+91rmIrb1481aM98ACNZUPoTyseaoroFLkbHpvw5oEehNaIiZ
xqpm8cFDINHSigUTvTn04gBNW4xyPYqv1lBCI4bjDSSkOz8WzDd9EBasH59X2G/zxK3WV9ESRqB8
BmdCfLEL3A/Ah/raWNZ+i2tuDL6OQ91za1qjlrS4FDajWHw+uZHjHRYsQEtAEy9c99Fxb5se6AuB
HXIOPxJR5OtpTDuvZKHGhQ7v7oy/8nwQoD3y0zYy1dv+ifxZ5Mh8Pk24I7rdNz5WRC6gddY2uvCu
6zn5Zv11zA0qfcxZT/cvMlfO5TXtzJ8BTCO2baDX15wgtReBqc8kf+Zfhs0qmPDgXClbIWAhKUsK
mWGBMGJbRqh9umPRj9HjIjmExs6BF6FXEh3FLoM85o8FYPCihTCS8m5tH1ji404iaHwYbdWRSaWr
KnjPsDDiVBtA4wPMwucaqIfT6htqnViVPO48lwMaotpS/hbK5ouW8ik9rFD+wdThFx9tVKvS+JfC
S/9GzKW2/xuRlC9lEoCNixYeBBhAPMBwfhp8qUJ+cOBgAJbhzIhh93RTrUB4raidDBe+HvNrJhIP
CTQD27V8TtFdp76hk2L3qWfypc+XdTosUBUltUHcecNaQZgvzX27w9bs6h262CRIO2q1f+hn+amS
UnezO11R5cgj2dEp+AYBjtTw6IUCJy8DPLxjsOWZQe0vSrTitp7x/foLmso01AV8RjjSLOTKaRxF
IgV241nXo3CkiV8InbLyd7RjfHugxnZ7ZOp+huRg02cQ3/iYI+wsUR2TsHrcLsmdWO3awHRaEOjy
KCdUdG1waOz8aw9+CiCFdnR05ocKDewBL60WoksFTrWHV9Aq8TPsAUJfdwgYxbuoyUOu7EYn+iQi
eT2E6lTag6ywyZ+YfIGNhkqaZeTQ+jMKimAxBVuKSVEi2Z1E27ksGSKkNoQluZv+uuAziOWulPy9
aTT8DQ==
`protect end_protected
