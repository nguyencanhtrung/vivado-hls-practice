`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HKktfuRXNLUhr7k0fi50JfnFXdL2vEAX/nsClluRHE4CrThVgLeb+IzojDDVFDrhuAhSLLNpg8JD
ALTL0VQWwg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N5Rr1FDKG83ZPdwhZbcAEbVDVH6nOILKblj3oq8ZtK8+As0Se/A6iMSsuXttt3xFVGqSMBS7dvG/
kusL/8J0P2SXQVaC0rNrpSKYp8RErdvVLfqjrH25mYOsF4sRKIOyN8LBOWgeRPQF7OgZb1SThCSC
9oNwC0cd/TDy5x23DFQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o91OoHW6u3GhhotAeMsIyLuG7OF2oIGI1tfJYcfO+pxRVIiWnmBgpMJSUoT3KpgEPGLhJnyRSP/Z
enBDX3cmGnmemljPQzkiVCMl7r1GSzf/clytbS0Aq6V4UK+u57MX7K//SCOQaMhaD/+/SVXDCWB3
CfPWF0gg2GCqaQbTsc5GYZWkazOgaRvUCybNDrMYmTbbfbVOle+JEBkCUtwxz6p0mLZzTLZoZh6m
jjzs77l5Zce5IXSQzknGHNr9wqE/RBsviBPdkbhBG8jTkTgScCHy7UsCEiJSdaeRtpb2+SRA87qa
N5k8SmsDHDRFPnMtw2OKKvzDt0Ys9zoDaKITfw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YxNF7aDY95YvelJMyT1cubgTv4G1i8H6fzKEb1O62Lnew1e+r/+OSJ0wCsmmfsLGjY/TyT6cU1OU
uoHYWGA026nqBNb4IckE3EUa9+wPndKfTYc1Idv4/NjmgbnBAAWM/d0gaqh+MmyjSJzanfmyzIvO
CP2rbPOZRuEQx+9C8r0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pfkBNOmtocxz5+b+Dh+IqwxDLBsGdcSG1fpga7Ms0atb3sKOLY2tx3FxNbT+yYrSzpspFlxV6tIp
0TsbvP1y8T+uJk4qyCfZI0IJcUicqqEMZ3fJIG5YcHT5Q9jbKQTP+7TQH6PGFyQaNp0xnjy8Cng+
47IPwW56Wr9ikIV3tM5PCvIuzR3mWfj8seqmh/nd10auIVoD1k6nNW+XwiSPjXoODKPOEuILnkTd
/2b7fob0jiO/5vfi9J5fWHV0wL/uTE+sR2oQOOBrc1bIuoKj8ns8O90oiddDTOwV6wxAVWqTNm7+
T7Cmd8/VDfHexH/SFK2KInVs3Mbm5Ip4hM3Pmw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Xgvx6IKYd9h2VW7lxk5Cz5VOGyP/QSST+2VNUfO1UIrs53GKC4sLxF3zt/nIBQ6FdZCIBDy1a93i
cxrEe97PZ27mtibuX0Y+uoAKM+uDQO4FUBdNpAr6S0vyFJT4JiUib81N7MCj1xTtYddOlVBNUo8M
Mr8eUn4ERtNLkZZwSFWfbdouhVechEOOBuVUp/vMl4olgYvnyiHx145GwwrMmsW5RltHWvdzJR9Q
PtbA0ru9/sr/DhSIkMOIZ6eMeiTyhzU3//NmoxWT1epf48r6wx5il6+OXXa2U4UB9rTfkyV+KHBa
AvRxEiMVB7AuvejGvyc6zlUiG30D5K2PToG8jw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22080)
`protect data_block
Mr4vC1z3vlqM9YiICsQry0ktE234OWPsmfhwfzv2xVsg7p5Z0T50BTTatE/p5+/JHXgxIX3SNTpD
Srp0vqvuxAYrtfShsJgZSaYfh8YlmMl5rvfdCn2xe0hpSSRcOLMS8dUbnCXQp4kLeys2Qz81mJ9o
R10pDAmS4a57XhQqY/vIYNiAAZih56HMHM1V8taFUAvuUSYan4eHC5zgla96wIGxPueiB/fEapww
LLO1sadDWB6bszV7U3YdbVjSqRpPsz10zqijIxT+eOREJsGqOlhleHlMRwN0/22q6K7tB1MkcNqF
5fHD0fj8VmjlrHwUFOmoaAJdfyHLFOTOKY8lIQA/hQC3ddFtPk+5lD03MjjjiZrNVDwrMbM6XGVC
VUwrTOBLxV1loh/OeYrekIYVf4qwNIKpffXVnFY1+4eoUN+jQswMRjoVrMWcraoGj5DzttP+Mr0W
dFgrRuEEEvX6Cn0ecMlgfd8CDT9LEMSsDff/N2BtabjrrUsfWRgKyE6srtnewEeL8igNH2j8+9qu
WRHhoyzSjcRwuIhqA6xyeMxB3wcg7jQcCOzdnw2p+GK77T/F3qgMMpCT7xc1p+maMq1H/9Fo7YNq
3R+WVxF58iAzzJncoQjjetVmXvvaMhYPRNi7W/8F7KjMZEgJha6ScNlXe/O9aOXSenWpPKY4YELF
s84jWzzrLqUOtZ1D8pjizBRamCQTG6dTzUeGJm7GrTTd6crf7X7o/ZEw6XBiXYfbwGxKTVzjkGKK
AQKjQiLdaIPPuKQbnlW4Wnh8lxPv8aSpAOLtY22JBGii/bdlz3/iydT6RIiOpvBhvpQZKIOSyNe9
30k64Tj2GULWrXmWD4MIYobeb7gCltt8jfGWGChOSbSMIb7o0s9RnQv0d9ooz8hhu30Couq+JtuE
kIeMU3XZFS+Uc/1eSEvrvYNAbdkAkiVQSzg6xFANWFAV7eM7iASdnSuVfavsGT7SZflHOYiZRweO
5KiCjxP2VVwSadTI0JrApAr90YLGJ3TQ8b2hindLhlDjHAp4lIRnfPk1GTs9oU8BcY7acz58rZee
oqRIbNnJI0rh3hb88x6Bst7C+Z0anAY6/Kb2oT5SVB0pLLJG9YWh6UWkK/O3SH3/ibm8yfs4GlkA
P8GdEtjCL8TqC4LRoIHJM+7m+DgPqeY299uBLYdFpqSnx9T4xs6iT+mq2zJ4zYAhcW7GkT6vlnYW
TkKQCEWEmcuahBI8PFl0c+XGKbnEqzJe/Dh1TVhXhaicxvspwo9KXJN0biGTGqty0TgAVgc1tiKU
lIFj0v8t3R4KEywYdHYM9cjpDTmZrH6ks6y7p+QdGqEKCAf7jUmdOUHsiSw2uylovpI0XBEbN9UY
9//n/xoOte6SvHUvsnM9R73doC/WnEWOAMOHBalu6/XUgUfWuh+//OXz/aR+2my+LX6QviYGVPd1
1zIp5wmnlWvZIITb/27XGkrKotsti8wvDg9smVZmKEe+7MOugyZ3O6UTQuXjh21dELGccutrGFQX
M4M2zUuJqwrZ34yksLAZ/nt0zIWbHx5Z3AZ0gnLsaIbVd58BekkInAaKi4SWpPI/FkQb8K/7kHnr
O4irj1JFZqamLllNVPYW9A8n7uRv6yb8tiKRAsqynOoh/gA1IiyGp4OogQGFKR3ut2poWA0m26Li
hXcyy35B9acBz6lLHR6nr48vfLyrBVOi9FdxjkDarmxoMrYasC69ESbTdUoMoZKMtolTYBLz4Xcn
AYBRw9G2Q6k4MBYWYFYl5MjkQvVi6ACgfneNo7qaMYfRsTNEXC65GT1LjIWKci7OBAovTGiioq1w
ztQIvn6RMOrS9G2SZHMzRT7kzi0rxdNAlzyW4lKwTt09PexdJ4Z6PRhCB/GrnrGRmPC1vC5CibMR
iRKXoDQk6rJWt/HdPrTBImBKEhZnp7kyHYvL88M27UDfXYWamrAebSDR9yIJBRpy4/8VcbwDjGpk
IHItk7kkmZv3e3XVDTGLmhLsPg1owVkheH2k4Ssq6LZ4h/Uy7XfrR0X/emuO5DHozAhQQ00iwyxL
DxfgRvybcIDUKrQkfXmbaEMDzUolME1+NUke1XjmrZ15Me0lGhRokQobe1bYcVBS/ZGuTqLe/+oC
HK2JplTKvZXPhEPsAlqxUBzvTwdhp6zYXOqCuooOHazDqgPkOq+KB2SzSf3VQ8r5iK4pYNjci/dF
Rdn46eTrCRvPcjX20sncv0yAAz8NaJI6Au6kSwadvLtiEnXDFVvE5KAj5QkYG0netrskzKkGc4u+
sHnjYK+ydbA5TrbSMN8jqijJd0cqrpLYc/8/YrW84nOfOmVzCBanbqimPba2A6HNbkxSBhKKe0jS
zurWcWrBmxM/zS7o7Gao8KWoY3G4HuJyUwUfx7muhRYg6gnQ9eIQx0inPZi0XsqCDuPVNad2dN7H
jMUv4H9rI/1nNghoOgZ9IZPnHaSCcmpFUjy6wPDel8UynCK3GeiD0K4bO4wAm8whYA46S+X58Ds6
2vsdnQORGkohw8riEgk9ykwt4QIxeTckrxO3OKJVWt6ejaI6ttcCLPkBYlVXTFASdUua5nQI0JV3
9ymcssc9uhy5asSkNaINvlCa33ZrCMS+JZiEBYY5KnFA0MR96XM1rtOPPtrZCbqRvqCyqxl1kO5c
YLHp6qsjPvRr0boXvk9gMcGQoqSD3Yv44ejK+FojlITNN4A40IjHcZ9AF1e10JNbfDgC3hIMZizN
T1H9paXsDBrLhvFdWw/JctAAJg8Q9B2veL3AQ0oewk/+60GWqodZhlrhIaBgiSJnUlhIUO6XejTA
1/sfxsj+Frc+NLWJmtLEEBF4TYdk1dOIhfklveXI4ef4NX9KxyCUAnpkClxpwiTbmG5v65K2ynY1
LmjtHlCcMYGyQOmJ5rbPNraOm/szBvHU4qlIDaru/VdZWfQt77HJsVdMBBHqZLZzQlPsgZkwuc+0
GeSL0ajRFKfdKqYvlA/1bbC5+eAeehcEm6IYJyU9Q3OLhM5dtQoorul0660oHF3xn/bJxEGtBpKt
R4H2lX/BKfGF5PYJ7EiXJnWD956xAZIDzHt3cW4yEaufI4stgOlOPYGsk285V5X6lGtmFmCokayh
8B5aqDbRkzm3O9ELnpTDWD7yHdxwneFx/o7OoS0mItQvAa+5J7YOe++NA/MH7g8YOmsQ6utYZLat
YZqXQcLVWB7Z6m4jdxWuyv/so67WFLCzcgVvOkjEHgUUzRhNWM17be6IBkXE5oHY1q12DEcqVPZy
IC4r4PC7+C2H6V+ib906/mSmyG2AgYyf7WAKu3y2FUBze7Cq7qz5do1mH+/C2yN3Y/hw7he0Q7md
Jm722bXsC42HrNOUif9K6C43Ite+omSMgJXgqAdettSB+97kJ0+5ML0z9JrkUt6DECiYfrBKTMHL
RZkl/hvvRIv7smyYZoUx6LsaQsBUX8E78tVDDVBd8GmcbOKdP2OW4YlsyCrvxH9Lnv9AYHS9zrDd
eC8y1wbRPhGMD8JACPWCXEZnkId7KtHkmtXvhCSJjFYKZI2XIHHl+zQLbQv2NQutjglH4XkOvwFr
ZdbFvnmcEU0/3TEPlDQozLqL9EyFcz8l0ORXKDo4Q5Mu3a/RYWy/Tx1WSJkQws9u1Kv3Hsv3rdrU
/eVsx0kMHuhRJIABKzuUKU1csz9ID8peoamyQxV0pg07PG4HZAVbmTDg3vtttXW1sLUPFjKbQ8wM
8fI8RJkq7cNqRG4LKBGeXe2XQ26GMKT6zw9uk7CQrP3btcggAi3hypw5aRqAU+NHLDcPpZaJb5SF
mqQMvpBsp9sJ0rr/eO1H2ZSCTZkIrPmopS+bVzMzRR+eQerBbXdsA7CEKWGNjUbu6l/MEe5IZ58X
NvbHCgxnJU/Ou6MXB/KkJpOD/S6pIKrXaETIVhSmgoD0md4NEi5VRtPNt8TG03alYCYc6R1pftmR
N0zByxyBWO2HfcRMzZLeEAHO011rVo+aC8K4QGrRvMmWABwQu5cXjdMMBiBWdWpfYkSv8bkj/ne2
NBZA+UDecOZJ4Thtk6HUs8w37UhPIMeBdFuiTEsZnz6G4XMJwiDWvwtfmrbzOmvG00hwZvpmSNht
tbiBDNwsxslhPbwq3MxgPR/1vkWf1nHbITkmnY1zcYY1tWLjwIATimlvCwbz61gn/5IgtOrFQ15k
L0oWtBVI1Es1gyRCpUIH4xV93iam+0VWjuOkwqQcNCx5tCNsbYMg89nWxhyNgvnwWPnwU+Ph+wI8
C4NcOs1ZzgTBOlqNNC+fv0hPIq5jtWlfnrtVfO6CPPwGyu7gFUYQgyRIqqsmExxsf1uQ59cx9clo
J2LwBXrRrSZVA9v0siKGSdPRagXt++X6dIRWYndknHmpg/MCdeKf4O2i4SeSAx3bLndmmoSDrKOE
1MZpdH3Hy9oc+x2YmPeNUZ1ltsjcps2u6LpvB6BOMqNb82yCLFekDXcaKr7fQ8EJs5qm3l649gIe
57idV8iuusXtgyKP5iNYivE8hTA7w8xeUfW36o+3BpQwntQL32GgVFgHI5zRaa4/9iZTTlmfYgf4
we9m44C6T9Os4qiJAENijkWQkC7kTbbJecQ9pqqs7Tehfos9CMCgIkN+HikCL6oTYvOug2pYGzNW
WyL8xcU51yySkUF4PDO1x4UR76E0ifJN5e49jxBxUflyiF+kKPmK4sq8jW7tgUTbvt410/ulbtoC
urQWhWDWLZ0URaqsBcoxss5o4rJeGcD3/f/qZIXNHHdgdpsbuwpCeLxErNJHabT0GdbYf6ZnUwyw
kVnORr1oe13S703cnodX839iKsXiDN1tVMv7+EpVlXAkJHSKZcRXNb2rNKzQW82vUrnuMTTKSoGd
3qamvptEREPIwFzsO6NBnOuP3Jj8qo2akUNw/texIFqABzgflvg0AwXEjSo38kAbIJww9J5GH+cP
kF046dzPU4d+U9ZK+MsoY9AgxJ5eRdMovm4D2gcpZqQOi/sr9EO7Fj74MGwN+DNPIRdPCG3qvkxL
UQBIBvKYfNRQsSAHHVJF1JBBr59cCHEJbJZlzP3oTdhOJH3eM1Bi0USOqPb7+nprsxQN8Ii/x8WC
uWgp8XcfpSJmlFqPYxCumkjRdL40Vwuj43GnwNdxzFhPQ+WfYZRj+IKgk8LqvxeyLw9GZ+2WxD0G
LpoD0fJbl32Ju9gyVIHfl+z+Cgz05P/zqU1Q8ou6uxxw3Stok8YekK3ljhSLDbf1bKE72BaYPGKl
7VzBAZiZW+axsxHLuAJf34xGx8JbCTdqB6MGQRl8IF2rsxRchr1VeLypc22QPREIzzyr0/LeomJs
w4ce+LZBGroNPuo5RCXVwF+BSjl0Degh0+W7fRTrRSBZw0XcJXN/O6ISwSfCO5wLj0541Wz2X8XX
f6Jisg5u3uG3WqilVYKKmNRINMLm6AqJ3kkwegC4qo5iOlIHNWIJqErPY+esaL6SyDnM6I7s7VJ3
anOdj5EOfpl3iQ96F+eS0+Vych/Fa2zeMmHZhtyp1vcZyS0kYl6dhBL/zCJ4YwQCuo5JDeDIo9KQ
SrhUSRdNdvF5f8qThRTqmkvtqFLtrM0e8ngYMFUDBz3X87XoyFMPQMNL8cdUmS+bPxgtLmLjK2vT
aXUatKYzjzc7InKL86R2UNpD9Nkp8vCAtvdiFaPvic+We5WfeSrORkLWvcFFlBdRGEP5nE5cjZ9H
mpB+emr9Oq/NvsS4GM1ppIxi7dAFDgCc1j35TMcfdWNhSLBXXsbF7DlnHf1bZRVZIjhn3V8oF9CY
bqAFIlstdPIiHSgM9h3gsDaHSvu4qSanM3iZhX0ffOGN8A1yhWgUzA/WqKXyQcDePfDOk6Y12v4p
veUBZW84jYGCGG5snqyrDJoD3+LPVQ8QU8xzyKr3OAGKWzjL2gmBp3t2dBQfdLKkSerCDibSbOKB
QiLD+btzuZ2soglFhPYuEO21O47LCri8CxYo9+0v6NB8UN0U2X5M/Fqe07PPPBhdZ1H2baPfCh8L
lKp4Ek+PPnmilhfnS+N0Qyl2hwQHOgo8AviyvEbpKwBfAu4ExPJ7TwEgfXAbjloFdoW3ygD3ofc2
XtR191QzX/ttaQAjKMlkvlG7/sVxeW1x3qi8gfBbHE3QkffjzYYrP7BU1WEQa949CsvOg1AqRxEb
fJZoAbN1/O613ZqEMgCtvLEE1x4ypzwHfSlowSHQtApYBBtVFIocKzXNg+juEDC5b++4eUeB0bCG
OVro9dEQuKd0WRFxYCIO/oxUUjpYVSZod/cI2JS3GCEHk6zMgMPQ4IAarY0Wtcbg4ffPdPdZ2s/5
WNYXw8KnmCXEdZWBGahWQWr45zElbdt78rNek/BGEVDvcHSZD/F34JpMuY1NGGqDUetrvpyMXAB0
2IAR/8Cesbcc3Yky+G77S5Ego0CpVEXIF6iH9ip8UdNOu3Hx97WdyADlOrC6P1oW3WWFIylmwI99
5W1drDgV5p5YuPnvfBLyNBsaJG1/LdTn2jm6oTFFrDwCLN6fuuT1WTABoDEt4lc2f2uOO2irrDn1
8wfC+l0rK0J3CpeVVnnl4fMAITxCsxhqFMx7MZseVaMLuHyO3mPB050oQCyAk8svOXRIoBCtA/od
vDq7AR9eeukP6wBdGXj3fnblKtyAEtBr42Et5kK/G1eDoAbF+W0w5A+lBqLbNRv8CkmgsG/YIyF6
bQmT0isr6v/JRd51bvpkbJIK8B8X3vbqWwqdTRHkZmesj6ZRKoCREF38SY3sPUqfW5cSLftsTc+X
0mwK3sSFy0KomXF8sfw22qPFiIgQP+/ZJXEElhc/gT+wuzlBNfrSMfDhRMkxJWG/GADNr5XPsxaO
ILctFVHNEoMQwRdDHTGlP1azYkseCkhkEzw5I33hoft+vQZbf/kWvuYIRrooFWk62pT2DbtxJ+b6
hGf9Hc7/MY1c5rTYACOw18SKBDP2jFHzmTic1rGlXX/KatRPDgQuZf2WrjdUaQjXgXjmbQkbOK0D
pYa22D5ml9Ep1dgkBfiIGTGvKiPILboTkZ+2zDdT+Bu42AQCCHqXqJXySjAg8kHRgRTP2zctNGPh
hC653it5h5J/oR+xIYzaGz2cfTowUHy/pbD7HgI65ZggtCrw6zDSpvWf1AjcmHaZHM0WMmi95MCt
Ijw8LMljsPfYLljya3ydT4k1dEgMrnH0wXEGS+I4bu9rvi+B4EK4gow+r/GpIoS6y+Sj+R9Zx/0z
m5T0izjHzeRfKs3farLEMT6fa3SCPruIiL954g38EmKg1Dstf7tOjIteQiukb97/L9UpKS8bx5WY
HTO4Txu7cpY53Jh1e93Yxmi65CqW/2z+SoRED1ndA7VzwdN5xor9qzFmhRr5c4QcM5xLZoY7G7EX
MlPQxH6wvQz0TpdchoMN5dNzu81s7q9fz2Nf7Xnipw9B5IouGaD0DNBdoESx3g/pqRIRe9JiFfI7
BGvyMhsWwNlbBECszh5+053Zj0dYX8nsTyE+jSUY2p2TIPMcxzc52J4+2aCVHEmXgTwyIIaP2KV0
5lP82TMDbYqj64vD/t8X3PnLOJ/TZLrePtzmEDWyNydBYgT/3yNMQEsoSxPWr8RQRbS9i9tXRcu5
Bw2g2ngqr/WxzlBu9sS7tgIRPiYS91FF5bIpfZGnLPiHR8WABdwVUc/4eW310PcduA3TN7TK5U9e
tfmFjnquQZ4OcVmlu/CyDispM6gJTeSxaPR0fPgjV5qEXtpbHiAeoOXnRFytnVh+wSXJRMtMqfm8
jQltRwuUqBYTGUS1ApYnzMPQmCjhjajtC0YEFBwYtyYXPlRw52EXMySG4cjqbs1DAdS9Pi5o3MJe
FxMcIKh3P6lUfu+Qv/URqTova/1xhz3s4ZoUCJtQoN2F0UuVHqjd2GnjChNvvbROUX7X/JEvA+qi
bm1TUjmowtAiZdwSTE8o+SjbF+3kyCtXPrjbnjus9o03kUjnRYwqofMyhv9TUVBfmFZBjH6ReQH+
qjoRo44Nt6QsQRWIUkjuQt75JKAWOqKvflSLcyQnHpghpJWlK2P7UaeFfxjJ15zP7qKLOglfLi8O
NvaY+UALvhNib40EuyrrSeyXvyu2qpQsqIZ2GyYfXXwtIXYVZnqNzrTxDIFe3WHG1FriR2EArYZL
i4XTw7ibV/z+iwTIjdCEQ7PBfOh43YWrnXBOMc6NXu5WIy0G4fOyiwhpEaj4vDd13qhT/C9oAzqR
mNhc66x04Pxgx+QCgglXN+2B9KIoGPa28+O0Pxh3VEzdhXS/9VjtXA0jjQPTa0vIbaUcj25rZ6y1
YqQRYeKcKSDZmXDdJV/NPzBRmlK3mboK7AQkOrENtfSjZX6BKwig82aMPM7HNQpoSOPFIq0Hboqc
kHwK/BCgM2jGlclpMcI7lNcc88XSDPLW4kFJilWW9M4YTMz/hqs6luaRgMNetnBFQ8Kth42MDVA2
4z5N8XViimd4v+BbOpVBL/6U4iQ4oxD4eIgZu+e9uPrxDHYqnCuIMkKYr+jNa6MbTqtxQGGSOIkh
5fj5Y7K3Vr76QWt79Z8VgJ+9gpeYLnzpFUDMjBtzprblFZEoFre2mj7KdAZSuL3xDo9StZ4PX6u1
TKYFff6Z2d262Za/+S9ItzQILX/SyBt9XPOOTHNydQ0etruDtr9j8NyL5h4UQGnkJuffjt1TG3nR
F6Wb+rfrnJqjImmk4Cyx6i9LSnI3y8dmVEzjfwBv1oquZtUsTMxTpVYKtHfohBeb721FIZCRIWLa
az1I00tq4GQiPH4O2yZDgddarSUvsPegMChXcnimpfrpHKPryaJ+CjKs/HhaMTuDss4SLbqBOAur
eS6dBv0X5jO/jhvYYPf90bAvr2nB1vjJrTMO2msXkHF2HKSIYKWj6ZWENmhN7VrU0JOBnzLdMCEi
ZGMjkNcppukddO1M7H/RHUhXh4YMCrrgu4FnxoWsKRT5eVp7sxuWCRWkoBoT4B5pCBbcVoxzfk2n
mPwJI/96haA0QhoLPxkiJLq+9w2XuKEWhKm4uVRDeAn/z5EIYwyPHj+4ZFxCt5EZ6aL8b5VtUF0j
7XoNDp0NA+GKJ1V1ZDCvSxv99cfRHelfo9zHVmAWPkfzBOHT8mp0ILfC9XBQgUYj/WxapO06lUOU
BIvMW2Zv/si3yiPWVARyR/X+Gw1r/+WfN5HQlJ/0WuDfQ5HIs9bpzwZ8Q67DIEcU9bTroMyjYtp1
qttIPxHHFbWU/nKj4KfOhzB/j9ZmPBWX4qOzD2odxiFF1bEGsGusqm+l/2PAGThAf0Pw+kMDm9LT
vbwZmEWBw+MdZpn1LCxeWOHojpRULJm3Wq3V/6jJ1WbLGKJH/qwLmAx1O4bV6Cm4DB/o/cgYlGIr
yP6i2bTJLjt9/yDXA8/FWsSJjlThwRHOi6uyzFlHZ+Y88S6p93w4/ZCXC9sAcPjBmdMfOgQFRJTK
44zMI4R5A/TXl/33gFV1vycBxdn+FFzeH0oBS+Jry96EuJjTQ9icLAnUzgEN0jrCevBX8SIMPclQ
lbCrK5W2wmb0c3fQp7G6ik5e/ZnhLZYv/lZLWoCII7auLYsH4f+VBKkeQ3UwuXecnEIwV8Kpa4fS
QkmG3yGpJsPB0LTHCdCTssVdy4Ss/QJnFBOjxUoySigJ4YKF4Co2mOUdrO0M2N7U+nfxQJNgtPlC
a8YkVbFUQ44rsf6P18z9I+Nzzh7jGIohtJ/Ht+ASMs09Oxsr7kFutWVHd4udyDtp7KQ4ip0rzY4L
Bi3Ba/ndNgBRlGibNPkGacQZmb3X6Heqv0S/iuF5yDYnLu6qpzqyKtN3O1u37Ucrieez2RoxrsKO
JCFiHiQ8QpqnGlnDuRtaijB7X9fRvbMRdM8eKmKXu6mHTHKe2HselbzEpyQ/PJOQTIThe+z8dEy+
UTWnBH61MsbLWzlcsd/awuBShzxLsaTDV+fcDMtAnOQpAchrhxpry1z7t75kKaOujC4yp44c+SeO
K4Y1vv2gHoRJOPTyOeTZW8cXTOmGP97MhzwctVxba+YMr2QhwYSOARpccdneIeOVwioIeg51vRec
IScw7pDv/43NMqebff5EKzOm/n/K2ew7S3AHk/7Bblkz4ISwht3JuQ50iQUDZu2khPZKhzfO01wU
YbZ8RRY/5j0bi8SVR3tqEKTSw4/kknsAi0Is0mVgxW7AqBAcRNCHnduuXoC966RaJPKbrxBbJf/w
DQ41qhUuav8qj52vIG56XfJ/KrMVvBsGL3t6Vi2iPiPDp0zQ69L5LLLFwRw5zYjBShupL0RkTIKG
lkCbu7TL9ijBf8yl3Eq2VIz9MjQg/Iz4Ix/oDh08uFB7AP1YKAQNwALpJKk+sy/ulVG+Zwkwujyf
y6IynXXxui2MpdJjeNV2QpemP8o4xFVLbI00L1U+vIcBQx6Ts+JE4lyrt7xuR4Qf8jea6NvyPohJ
gCOinmYq3hRDIArxT6gOr4HQGkpLMim990eq/Tnn+8QB48PRgBANbleY29NZL4119gDS/WSH/kX5
z+zO3eGl+13Zsg9/ptVtAXHLX5aMMUzW4Swj/8SlnPi8yHWahIwPPNLuAjn7PcnoCImSmnGQidmc
g0oh+8bJB6GqjGSwgtt8AmhcOb+Hn2aGgyDH/sIta98pj3z2tURk4EkMoSNPqQAIB1kGRa9CCv7m
AHpCQOsU2CZZ6rVsDRlwpdJDm5FR+f9MJNKmaFo52BblSL/5KIehT84TEzfIIbrdl6AtKNIc20hw
He7Rnjc9GnL0TrUjkW4wQwuVlPK3WC5xxPZ9TKjTbl0WyXC0sHphTtKNym+0Djq5hNWkoTY2wKEe
lUROBynfGW+TYQ79ZQ8FuY5SNUSghIJ16mowGEag0W7WIe2Wb8zb2IME1KVwav6rer21sbdPEwSQ
+DzyYllN6JqFZXTaqaLp4T4GznJgVJk981FhkVm4WiCcAL42jlewLEqBbZkcgw2p17v9q2txCXvq
L/j4O5YzPejEP+0Q7Qroxz2Qgdl6MmGI/1bKoFPt1DV15qSw57DQjTT5KmZiemNBESYdkKfJ1PdH
2WRZVk8C9puFDSwhzAKC64XU82qzJ5E67srUa8hx8K1jhZ6u/6KDOzX0EBlJZcuHyZ0D+0j9WPn1
r2Hev/ywm7nkxf6UYzVmAbfff/+Y6W7Zvq9u+5H8NKwb4aoT683Dy7QpMbcd1ENU1Sp2mB+720k0
l/1scLAT42iMLXNwyknjxKZHXjXTcgbqOO2kAN/shmr/1P4hjrlGswzfWlBS9VAuiOyTV1rvLOpJ
SmlD/8+mAo5AHDf1zVokE0oODmQRXEk9UNYNypy5bb7Mo99mF8myZ3txQk2YQeZPFVpm7AWFGjHK
9E2TrGaL0gpDe7m9DJM/V/crXe5zVxQpfTja0eTyzcwQj/nGsm7Xar8z97LVV9bnb9+kK3WXnzxZ
cfrdmtbp9k+NgVCtsARWT0ZOUo9QKSDQoOk5eksiu1ZrpUzy+n8TvlXdcMtI5sqSBjIkUFyz/mDk
v55J8+sxPBRKfY+JEzGCKqk1hni1otUMeieFX1sXWhwQNJ6rbb0GLlbYv42Pg0WTny9VTVKtEXCP
7cxfayTGQwAPPaWp6RFJa34sFMO99WwveDUwdn+/APtRzPDMhs3r2pkk6p01vUVoJc7U++usMffc
Xzi1UVoVejhlWCgwdbs9zGbw65Ys9LqMMPTnuxCnAdDFGFpQ7kcQdvXPpeBEx+EyIP4X6HUX5NPX
ubdJwHTheyAVK7vBbcieZNkk0wJ9HdsUkkl4vG1dj5Ap3amPUPdD8GyhmwHzDGcTm0gqE3HWw0qp
VFUmsfF1jlwMRuEXzz1Ws1E/9w+Tg/ETwDrzFqA3HyxXWhKD5IJn2YKbrK5iihM/vY+SGuAbSHCy
JKg1Z8slZWp54Ts6ZTJLe0ibGzRZil0jRuye04dW9xADPS0zA5NGLaLAPfVNgReHWM3rt2q7ATzw
g3giFz3p9b2b2USglrM062+ASkxJRHMr7R2jqN9JYPSFG8gKagcMvTbO67IKuGjlm5WdfqnQmxig
0M5ToUpWAbksABavRE5bLjnqjyJ/kPAKzsBPQJ+tRBhvLPK7xTavl9FkB+szPZzq4q/TiVBXpAsX
54uXZZli0akpSILZinyHsWh8bJc74822fumirBFvU424k1w6PWbaj0RGoFPUxCA5FpaM19oQ31FT
HZMlERZnULiPtPe6f8Z7uxY/rCzTE/ZGVGqoqv/cZ888v9EzfsQkq7zH/vvDAeN/XFewzHvrbh7I
EvypNL9Jgj9uGjyIGrkDQlNlmKBzuqg1U7zXd6fPt0kQaSFC0MzUq/6HI441otuWH7R8BU1B6/yd
WGyBNCYCh36YGO4HTJTZjgzoqRGdfaJiw7aG3WTpab4v05shBk+kN5iVrgo/AAczi4hRy9CQh5rI
UQIjeRuPR7r4mfNgKnX9sa42U0hLmD3jYaywyZrvnC9iiF80DlPWOUgZDe8rjebhw0AUPcJbaAvd
MwueALveEpqbF2gMV3dXSVz80wzh//JSNubSQoROizHAIxhxfjPORSE1qb5S3VIeoNqciiIxxSAK
T3oBwM7YgK2qjRNZm0GU6v5d8LluT2i2DEi499QwevQW0yDOg5PtROOBs/S6mlBOWIpLxzt05WLl
3rO7zm82IFfjC4zy5WJG2bdWzx+tgxcdSXKdusbVLI/J+2sWD4ls9Zn3mV64kshTcdBJphoXqBni
jk3c/Q12KhQSU31Q7rUOAiimQ0/fHc4U75eZ+DzvmkC+D6pOBRCOr/iRDq2NztIibM8PStXCpVvI
Wpok1HfqhwK+Wjq8SqgvYVBpbKXWPZ3M/a9bMzgwr9+LsGPbA8ry5I6jw0ui9AGQ6xp/2lVqcf7m
jryGMtQo8NQucoIC06rZsNkgOMOHvqPKOL03m4lkR3Q1Fdzx+EI+dDuZq9vthan0zQFuxt95KT33
3qHCJjhnXkqRzaMDRvDoFNBHsHZnvPXzzCdMuqGvJgWCxeEUw/JvJjEMMmv5mIcZXnJ2wLoW6LVZ
qIOVBw5cAAZ/Oil5zJy7NLe1DYQmfAzQyZ16ds9fQnEaoj/4YH8bZWQ198XvfSsn23Nh3hpm4Wag
sqZV4Bybk7iP3Kcsdg7XF7Z+dw2bdUMmEcnO41YWgHe28crn4NVL9u6PxKvzst32Ujnk81cMIaqv
LImz7QQWw0jHgSW3sMsxjzMO08kREnN1v0PB+dQlbzhtHyRz4gyoPiwS7jw2YGyYV/wrbSurojaG
LgXk5r9ltHtMc7/df8ZUq0n5rJWHCF+X20jLqMx3xf5nksVKZ0MdYWi32iHRKszGliCJvbNd9CYq
Fv18mnVPTrAJzk3lhi/W/AysyS/0N1IJU/bbZwi+uZeYU2MDelfNcKH00+W23p2EHqNdyk+QR9KL
20Ivkv3MxHKvTR1IutGkEg25HTYmYh6C0KwDKpT6McCBK5rcuwaojeTLUT0lL8CrUKaHCrTJqUI5
VESjIibWyra3nWeJeewN3cBdp6JLbFg0taiNc244HiD3WajXnPcb/BrKEo8BgFpbP1sgR57gzj8Z
/F5FGkY7Qf51tAcJ+nyYqKxr4+yhzDd5AVjOpr3jOXtw+drhnXNV7z9Uwa3Ih7yTyp9lZAcmwH3P
ioTS+8bknQn2PPY5npVm+/wQOaCKb3lKD73oGz/Jcjd4y29TKiHCrr0KpO6x+h42UhjL8DshNrzg
67DFWkiAi3TlFJuHq12zmgwEfy0CJcFPppixXIedzaKdEVGl4jQklXWomzBeqlhUrUykamvyNagi
FPMlI824K04RoPs3TpzNpUpNinn69ZM1MtEjmkjEDTuHwuNcpYK4IstS2vCRFGs9mxGdvdzo/ogu
x8QHi3dvbM9h57hqqpLfME6fx63PnnUfZtinc897DQtYckdsZx56pKITkt2O0JnRCmgfNoj1MIYu
E7vpIxItLGMxPmb4KTkGHgj4Lvlktw3kVf24TN09IRntVV2TIc91M2hxraV9YHkGSPyflnaPJpc/
Rbc/+thLy8AOLzy3+pTyReL2pu/BVPlYMvN2DeTQyYxnvlZuN1SjJB7Ha6nNrftzBo1YKK5viFW7
rEIwFksb8AJ+yOVUYx5XRSHouJrWZ89yibNoy1M0MAqx44/urr0LD6IZs9O+kBB53MAZbnXNt3lE
6sge0ssnqgAWOcRkFJqx1MoI6REtU2wUxruOVEFwsSK8Xnh57ovekVwKDyPdOsapOPYS1FmU+yB9
mEsiFWziiQ04VQCDmvxVZRp/C3zpMjmFNIsMgi5jPgJWUk6VAAIIy4drJGH5FVcKv9EICAB0O5gO
FTX8lcmvAPgwdLkUMOXxPNsTuACz2EMIqOfYFzQG/Daj2PO/4gC1yQuRG1muKAi2aq+o2Y8bLFWT
lHPnfhJ6ShR+eI0thzJH/fwaj7LdT4WBwTXbK0S4bbeYYTk6QQXqZsc+PIWnWcVIMq/hZUgTkVzq
e0k2O2BOymL+YKLaVNSEHHX3/8rxUXJeRVHbufFsZ1hh8xWWcawA32B/ZS6IwBeAGocrlrqeuFob
x2R2F9XoTbgWXbV9nZ2CFRCQk0YeLS+OlJGOIivvLLYqPsD+MWxgHqt83vRJzv6x4NWOsYuF4vOn
KkualRBIUqnYTJgjxwd9KSJDoTcpeME0bnf4gFGHkwLHP4G0PDOBy3ITQxcjVL8Z32NJm+MyOoZi
6IwruT2N4wh0GFmavpcd0udoBAxNKtjImv4OU9LnnMtdJX+F8Sk/NfquRqilFuIYEGVkDiRN5roc
XoXJ5KdWKfX2e05RQWs0eJhU2aYSghK2ojTbFonBhIL82JRreULQxDpRt8Qu7QwCK/eILg7O84n3
O7JDnJrcwOuql3dS585QzPtR6N1BRI7hkH6QPsCsCbMJbF28tAz98smdAjbaongbP3qbCufOnyuv
UZlPdaMtdtGyzd40bPKoLVG5ve/5bcpdCuLazThh26o0D+5t6oGYawAxpiSacmHskl1Cs9Ksb50L
9q0sRUde7IR4HVeuqykmTs0XGoMcrEtEqOowQ8bM/Ga+vjQH+g47eCFrcGiBQ5WJyHBgvRu/hJup
sM50WBW9NXeWeJ/f1QY00epQXr+l3O5GDkXtPQ4IZlnPuVDyGAvcpLgRKnt1XdwGkBZo/Chjskj1
LY4ylsp11EKgekH5ujpAKiNsu5cozkP7qbT/zKNHYrrxQhwgYezSbNd+zs1dyCJKS4aS91EyTQUK
9vpeEoUmtBfGkccsOcQiU+6CAdtE1FY2mofFxk+13fnqGlEoc5/GU/l9gqUUI8wJSte2UuLw7lqb
AvJ/V1BDI+iKtEr5Wk0/wBUNboUG4Fsi/vJrZ0oEGbqONPZME78smRrl36Cm9CI4QQsLZiytfbdO
G2YnQrbx3E9KmaYluSl5tVq+rF/EjoFH1phCgadYCyT2ANhY9iLZPolfZwHQ6Y5jmFj/P6AHigEt
IAbworqLZtEeJWVTVb+JvvXg8CWUyBjZ4cis3frJ7X5CGYlrISkJIiiCf50GGeLLLYzqJxe7/CDV
WYc8A60cXXIBmfpl7gQkojtX3fQ36fesxRQ8v4FjnYGq8bm9UkXXf6YNLl3ccWmnJbGowZcM9aBs
JhWq4/bA0jYQ2H3RjgzQC643DuWXWuMvZu8+XYuz8smUPuRzyKON1k+y4nuXGrwKMCokPkAL1SZe
WUWcIw+kKhX8i1HjcrkdJZvUhfP8+ptNHUDn+SJxG2qu+DtJDWW7MUIdq+ZAjQC0/D1cNvRJwO12
+k/HHSUh4mppCJu0FJ6FZIhjHh39Nb6gm4o1oibGSql3iNdCFmUJUJlUf77i+EuRWg168BBvVr05
hDDY8hL7Msl+MnCNf3zt+hkF07H5s83/bsDJWeIHTDko7B3drZr2vHY3V8c2U/DzBxLkENQ2VijL
gbWEQzfCSol2rpU45hUSqnW/2kvXpudA/zNseN4SBjGmzX5Tr4t6kO7OVswvMqROOsX56IsVD1a0
tZOCHFRJswVsCk3UMEYJ4mdpK2TbkB+qNpj8Ib+XMU5sMDQAUfgKtE7AEm2AMXeA4NyOoRRbwRjn
cT03uJJ0tlm2+g7IZT0fkBgkV+yOBdv69VO57QX1D3FtUQOX7iYoSCpDqJsYWjcfVeg0cLw7VM37
9P/I0SXrQWkIkf9wIRszJgDAp+B86rxdN1DzA0mgHRJJTzs6StqEWQRXY6m1p8XdT1mJQ9VJH+05
B/2OTH4RQSvJyY6jay0o/pekt+Sr26zuPsP3JTWXz1sZe6fJWgjiOsOg0L3BPqulKzdFPBmzHhF0
pp3bw+INAzvhpxPijw1/djmJhXjMtYwUKBBxmUjAeuQ2gLjoRXjTo0ISc7e/XxIgQZu0YbIblZGA
77X3D4duAvaQgjJrB/PDqPX3qQwySceTlKPo0xTgzbpDphg209NNwjaK2Q7VaUh561mmtEnfmPXV
Rs8WX5qMYXw1Uj6jTUFxVFbsPVMoV03VkFlq4Y/GlI9DbnL7S1L9faQf29cEKI2K/SPeB1i0csuQ
YRyVa0nntW9LLw3yrgW13LRyf4e1FomKwLU/bIFd7gTu38TGGPpGCQ2PmMtO14bVoVqEFSDrQUxa
hgR5CmX4TNEkNbSwDxp7YM2XuVcTicNU+wO+E/dNSJLRHYsJUi+YbnsH2l5EXyM4OsQHUtsGz0si
XezMwY9/newod1FREVhSCwaZFbGOKUucDBqgGBc/Z420Ln3Aittx7LsLGL/cS33eKcShUbuy4LhJ
XzijCs1pG6tZbClSxF3m21O2nf2M1fNQfyt31KWs5Z2J6hpuD9lc9JPTqJil3+d76917cFgvxomU
tW4Jm1VGNtYQvPyErJTlEXiyj9b6fRyZxLQ8BoigHirEatbhFkunak9s5l7Zr4VhV6GU0cJJJHhV
UmJ1gEtX7RNMLXl8bc32UIlD+fMSRBlrvR4rdyiI5GhhXBlKlqX7WgYU605UbZizTxdNZwkHusGK
43EavgSyHTGTvvogWGdepK5rZdxdW4qXUo2+zION2iQLBDOa+tZaHDJ/CF5JRxetXGoQGOdWjuE4
vS9aADJ5eNE8ExyuGN5Bk15WUiEZywU9WJgc+j329eI6M8wPsxFVS3RjO/lIkXIpy37NPqbSk/5c
ufzMmzixYPZLBE4FsFkKYXaE6C+Sty7F6XhIfZRiUUU4IlwTOPdXbnwTCPwzBVy4Br51917THOy0
XVz8IEvS8pSzsrLe+gWnvOdXYvYynRMcHyzLcJ77up3PRMbUdEMMvcLBpqeRB6JrB6vs/aS4oK72
aLYyM1hqYNWWQvjGJtNe5y6zx+CQ/J6b6w825LZmmzA+xTNzyKe8Co83aAULjhYxjTo5j7+8VLxf
0om+40eJS9HwhMMD7yo1Kr4UCY5zegICvrT9fNe4+OtGFmij5WcwPBX9Ayjbs3oAf1i07daQ5FLU
gJe/ao5sFc0ZnpQ8FLEMQa7FuEwrzjJgfTrORYsXvmJyvKppxJkrvr+MFZeNClRw+D3U4oYN9NLA
ia5sJHbKdZ+GfuLFtb033O5SkeV2ndYzXIWeGdntUJVJhpJowk4kSpm1oqNbJoo8pQe7qS8BJDm1
pU/PmvyCFYIigcOscWS2xeUpqKtPvz2eqlKuz9cswA/QrSMN6uB0pXy090n0oBIFInLKjYoMqZOh
qpGyDSIAj0QLrw1e8yvpTldhIXZo6guTOJx4899SVMuL3WNHd7XoXX+dkDqu1cD9+SXydZVUhsPS
yBgbVdrUy/ryxyeV0xDpP0JBnnZMSXJlACUApBMEdSvM/Bs8ch3YsTAlXl7tVize5cG1BsUFxYkm
d2DIK/uFeAMEzp3n4xmJ330EVlMDjHSI/0v6o2fZ2+yEPkdoskeQU/GkwuFpCoLSpbwsk0fpEXTS
S4vmRkRTg+hlfhEG8KR+75voIn4X9VZ6NoW1xSnxKLTY+STEorg5Mk4J8nvlT2qG7R5S9KUBBiwg
dktTGmuhFLuaborXvHdi9eUyJts7Q5xu85Zg4AoFx5CAw0ltSNnmXng/bLqlJYfarn6a0EWuVzYO
1jZZe+GUyo3rQ6BoVbYK/GCpqtmMSU8SelnClhuLz9bxqkH7OxNZfTfkJZ0P0Yv2pLXFdDk2jtlr
o3ySljL/esaFgeWmgtMOpn9UJ8rvbO76a3YsgxsHDzcSzq/XyowKr3z+NfOWt7Ubmk/wk/xEhCxr
cgZQodyRrZQDU0QnGV95hDFE+1BI7dKPN6Zb3uB+3D6BlckR12gehWAaz4JXoZwYszzeWZLcOMh1
KaeSVuGK4dECS0UCByWeMMTNRTjXZDmD5MLgmeLXddZJitv8vyBm+eFO7xsOrhwjdtMUnv+sEwU9
2hcxk2pTtJEdOi6Y+I3uxUy9bI8iiXM29Ts/UxnB6hm5V5H65Pgntn4UdFR7T1jmGBWlhYgxTbLf
1M7ncdIlIWtjtSsbTDnbhP8CTU/PYmQFx5bD7ZpcrfvlgOg2wPzkIsxjr754iB+nVEPahGI/R63T
DfL94y6eHzydrvdjqqz3JH0/o8soe3TSxI/Lp1uOnPqhMU2xyzVegbpxA1PMOHKjnpYctZ/QGygL
JaP0gMD+kwVVjlZeYFY9aE4XDiAzEcePFrPA3T6wLf1s0VdPuqe7LlqnWqX905Ll/2uPwvLPU++v
5dW4LGvGD6+lPdosE6ZX/C+laOoROwZ0rOFIKMIuhzKAG52CmT/Rq6lpQ6BncoBc9rDb2jGzV2Sk
Cs7TPegx9oZMqaZ/z8ztWQKJiAhApJ+EQqLOLD6HbMmMa2l+LfiIIV8mtO6q2/pa/wP5/CrqJSE2
OkthSk/i4JTJGENT9MrgCYDbjtSZ17NjeMG6fL4n3gGsnPohVDn0P+607pev54UhAPlmQQAbd5qC
BjRn2lFd4iGar7T1AcDd8rgnwUaPYXIpfL06gTuTqVKSyTw4stOPEDJFSb5P1DGC3mAfTleHSm7S
128IwfmPpkNW9GfmW5JQrw41g49cXNJ7TZ0MVxC2rJpcARXkHBK4t+PuC5BgBIFOuTyTUggJdI4o
Le3dQp0UE2RNrEkz9TAJ+sgdtP6TSefCiKhYJ1Ruxbw1tvmB5Usbt8T8sL4TjkkRJbWb4fQ7gFsO
RGEHzVhVvuryWfkPrZOyiPfG5/XtfN21+110v3uPhtN9pTOT0ph0HIDggJ5iumQMonYsz9ppO7kC
Nt70NdXj3yFiVaedIIdGtEJgcupKMaXNhVszeompLFvg4mx3/J3KClLPKbTse00TaBqSmB5+UPYy
UueQzYI8Fa78stvYSvFZ5o/Hc6kbi856WGUX2l0a8yTGXAkKDOw6oU/N+lQ8aJ3FPPIG1N6K40Zs
S3R+Gj2cuaHiQN0sMh5UG60kkMcbEz62bjZKy9f6oZcPIRXKqinx5FOh+V5OO70P/TXWwLr7htYp
agysjRPAgLQi+3jt49NNu1mHcvh8W6F7kuM5CDhOmr/hwfrdZhsIuevfnsILPq99ZELV486t3qrX
a5BhZMqzfTxrtwewpUKYwDakeCtJ2BhBRxjZ9ALq89pOBdEht7VZFityJ2HHMuaDtKJccg10ME+1
Xpf5urDlaW0fbXayzKBBeyMt62IkemHpmsrhKiEDf+DzYJubm4el6zpE4MOXYUlxZPaNjOM/5UsY
0bZAml7NaPHGxpDMAAe+dyUN9VywaK9yZA+Ooc5oEdP6rlgPeZQOymIjeA2MIKOUfQlMa9O0e0ie
Axnb/5KucUzgHZBCy91hJFAUki1E2IM75SWgboQdtEkFaMtlGDvHyv5cQUAA+I09mytZJmWclh8P
mLv+P8f4Gi9QSJ82LgQxWzQ3xw9QBt+bETcWL3QfWgrtzfzv1YpZjprCTasBqdFoZIkzdcwtz4FH
MDgWTHhmTgI9UxHjJOQGOrVFDPDqokMbOfOtKrnRfXQzH7jhKEWsWdqgELToziq6tMxpFUWFF+MH
6xxnsUUpQCHSQrhfEO8Ip+AfyVTT9NKUj89KvRAqHmpjl+j4IzLZbN9vi690oIP4kmcfA8yztKCn
F6RlhQYWuqwOgVrW0lbc/13ccZAC1CAlXlw/sOAfXIiree9wbJhwI6K3dy+oGfEwX5arPv8VfoJ1
OUA8Ataf37OT8lez/qU1lelwi+aFhBeuO8d6kEMEF3Gsqtus06R9M/ipG2IwU3NjkF3MF2oAWL5l
JuC4fjBlfWMSdNxYxUVZUgie21LCn5Fao9AxeQAJ29+UDKH/FLhekfDuAj1Uxbwp0DLNSIbrTJSV
8vfVWcsYwRro3H8sUEWagAaocr41VRBziLSUdZ5Temgl67Wuj3FZFgehTr7gS9JiFNHqr/4ym/sR
H9cGOdHMl9/qoVeN9nGLFdZxkwAix5Iu7/zrQCOUWq/nOsVXQ21aID/P+QlF/tr6HOEdYrgWP8qs
rzi+Oc5qLk2hCRsyAcoUkyU4lEYWvBUOK/tjNYJt39aeiZF6YFBXU2PbpOEU1ua4dodj/0yytLEi
LYwlycyRZwkDVUfJST+6zRp3nEP4EWs44r4NA+vgOgP3aj6N51gck0aEMuwGiJVOPrCz392UcJss
E3SYnMRea3PHqsN5KRWZYMPNqaaaCJlXSb7ruwdGotfuVrk40uWcg0kLPI3rgAQhbpwyAzHZJiX5
3p/2j+u15uBbSB2gyx5TBvKozDe5WGrnHGL46MpDkq/9EyzobmAeEsdktAtw6Sjjz8uVC6x/IoXk
Oy0oDQPf+xqW4Un7dy869i8bBsypCnpLxYy4qaAds6x6CIm6gmf1UYjqtJ9ZkLpxgSv5SDis19PZ
8fpFUFL47b5nKTkAuQAn3pOQ7L02U+5eWYPG7HXOW1xBlxsaMqSdzlTsy2MvQVMGrwWBhzP26JJT
ABd/PAdw6BJDmg7iFtyGK/GIVWJQdVVbNJcieir6GjmiGfLmK9DBZiQ0urV4UPSXhqnQocAdWHYQ
J9O9AT7kMIlBBr1VyTW+fUqg6mupDpbareLuhjdZ3u+0Kl/TrO1YIV/phBEnp8EUNZ/tGEkcunjo
mDWmvuspi2rqQ8SBrB1ZGqGEPfl7m5UcAlTU2j4eVs3jWoud5i2qChtnwvVJlC9rNQk9+GOH4h5i
7qWF3/Pw6hbhMdadtgXqqbot3Dln1rbMO4qxLW4D/JNrWT4+MRq0PVEjFjGypVdMKI4o9NqaTSnn
T4cTmBiX7SaTVC4sEwwdKKPYuEInGcoE4SKBZ2zeAYXJcB53/TzK73nuZYALo1mofasz/CbPyWsj
B0rTPMwzZMsDhlVqBNyHvxtLq0Wm8MkMPwSVGYRPkZhZQaL08cHBn9aq2IWIGFFx5ZFKIcIKHt7+
T7gs26VHuzerUrJ/uKRP42i4YUM1cMSDDTRUpJwA4bbR3SIC2fEJzcv3QU0VbqTWdmKYLVYRQVEd
VTbiJIBsQweFpLLqx79hyMSZd8MR3ZkrdMyLXtr5VaUMFOOHOh5Ayf27lGU1hQ7wQyZNKpFYV3FY
1+XOFycbmLvwBvTInw6+BQ0Ju2ffLORCKDphH0folFcQXRyHy0JHWX7xLR1mTyqhlMEetoT0wWjR
6e63zE8bl1Se7/NGeEoMxLXZxnJxESExyq/nvBlHOF1bYDzsqY/aCEx0QFGbUyQvxYD5mS9TaX/5
/ripvCDu6oaw2aMfPMaKkJWKLqXs4NbbRbPM7yBkP4tAd5ufsdeIVOVVtXeuAuIcxQOyBpsBwoKl
E/XW6LLsCfex0R//282X0ORVuHtY9I4tMSnFShtvjjN3al5KZ3HRgVX9vbR7RC3e4AO0JfZvqEpN
jWQVq/kw8jGKGH3iIfyhLD7N9BLYXBrQyuocuX8IJSsxxoM9MgoOz3RRYfzxmIO6lSgLXSFb0BM3
YMaDgjbIDx38KLTFBi8S9tjAshRQYuK2AUe4y5nZNYv/J9sfpLB5uDG0qFOkJ4sTNli4KP2aEUpu
aBkCTP+sq2fRY8DCotB4E76BIjWL2MaEUCU4M+idRgApypqZM8MkyEezERNdm/GAEdah6gesQbEd
HQLBew6qnDT7gXG/B+6i3cVh74TIn5gjkcd5yA3CB9psgGfMLtbBFUZC1bteNcNrzky3OJKYH0ST
aPbQ002IY1Y8G1ImSmZvJHpDITFtAKPVdi0m+7XSN85IYW9QSJuEedF4XmeIOlpx4z/VmDcYXKk9
zqqKcIxQFfEaHHag9YPX8VAqLFUywF10ZbUq8X8pdUslnqZI8UgYv8aoWFaKaNXGufCha93G+jZX
zHp+1kdhCqnOQ2EEYajeIPy6/RJcQIUXnIHr8klsBD3gZ3aBV+ZmQBmzrYDM/8HHUVB6YlCDW4XX
mcF0J/XchOE6HzIuzeNkuUT8Jqf+ONZXI3YoBrZy8L+CDUD6MJzQGcGz6S6XsiEQ4ijP5BI4ux/D
pB9dGIl4G//qwy2yAQRgTOvc4+alJ46qyMONyr7SRyAxidCOygDlELu9IGGqMSLOrqoicilQcwNv
fZucuZqedfRt1Q7eUQGFR5Er7VlOM8CH8jtD7gruG6VDHJi3nMq+8GHVDEbpgO762N9BNJ43GaQG
7mwbmyg41iROlVp2mOVzHsK4W7tG7+VgunsGAaaxSl18o2GZ+t4kwshn5bL90DGUUwqxffSpD3vE
MgwMTG+ijT6H6+hlYuLN30SJkgLxbAw+W2S7ouFtxfYONYUzvU5uN4vNYfKZvaeqKn8xJByqVyDH
W87pQjZJE8FFEJmiCGTDNZEe8df+8wWBwMb48EjNqVg0x6Yvl1WE0WsvqdwNPpsBq61gfH+z7IMC
393ty9t8AQF0jYR29wfOihUP6H3iyyHuxwh5FjzazzKaZbgOJijszpBcQy5xll7gcJl9GI7blREN
nzqR8Tp2XSl5X/A6tjHSM5NtUS7sOzFQSpjDIsVHvV4To+Mygafm9UTvgEKIatfMPIO+7yc8opgf
m3DM3TY4gzXbkvECPv8wptMxgoCX4sB97Ad3RSY/fRkcjAkUA7E4mcfIPIHQ6qGweKl3mgiRr6Jr
yTv16UOt4RXLGP/dVj5IaX6UQwe0t4A5OALXc4DIXOosnMfnmhyIhzGIM2GBBODouUnS5ZYPK5Xf
yjnvij2mz/xajkwVDrk/PwA7daJ+TtLheM97pKqQs/+wDh5WWPnV6CJirMTXspSOxAxUQqdF57pK
Gsj7laHCZS+yh1zRSj9+IUjTaWHNk7arJZkvcl/KGkCA9P6wcrN3YGhHTwBi129p5l8sluY9N4Fi
G159nFB3gMU5k8Qfi2K2Qf6749BRIcbO+m91JJ6KH4iRAclMAYV00L+MbE+McWQhx3Q+xQnxud7w
fdSPX4bciUx7xbGazLpBAbTF7Y0vlAkkzJyL1pPNjdT5xBl+MNbw2KtG4i6MGkjyjcWBngGELMny
VxM4AaaaFC4L0fzuqQ9zZ6vlsN/CHYCCwbXZAGKJ4ibvB0YMQi51G5VyU/2v5hLOB5jVFxGn9oJS
nF3NHg2sRaZ+dP2FcxXcZAq4WnlyHrTgME/AZTM/i8XnstxP0gDgSzFonv1PIPzaBm5z9AE4WFVo
SO1xCMfEybb/U5MNdfTdCzaNAH4mVkBnjCRjApE6GtZmzIB2WBhooDjTn0iHGdtl9xNr2Y5/g/Io
aeOll0YpIb+8bNlXBNTYqgM/SVF7mQFlW92LCa4eY9OkjD2Vr6jAfJy4K4Q64zZLZoHohLV3CjvC
qvFwJ+hBfJtl+waqNmbUVxtDQi3QP1rd4ZAQOUvadii4o3tS3ZIWu9ZYqiq00+WapR8ReKA4hYTn
+EfT2OEsIMA4+jdybPCx3rsMRQ+V2oIIk3aRYpBGfI84CsEl8Qo/EI1/5JtOg+mOkElmhnM1U7Um
jBWjhmR9iVv7H/hdkYfFZojV55nAvd8SDup7TY10KoXDG2rz6T90a1yWRLvUnvOtcAJvKt2iNbXR
VuxIZuupLh2WlKBJz0hKDvSRZNJ0tX/GpNt8p9SgpeqxI0/Rizh+6eYae60PWsm0kBNdkMyeg7Ts
xUqGcRTmBQFIZAKpI5OeOsZ1CN0lzmEzwaSLsLtQzpLt6LkwyKx4F6Qvj2PJ0PovPvOZiLaHMoAO
Y50S2i9/nrmoFSDJCk4zrPQZogbWXzbN5usfHb2ZK1F+6TfV5R4ncUZiOrD1QrJdLY2g1qWBxvZP
Z9YQnc+Gki7/oUmYZ07C8cx1lY065crHNrbIUQYFKcHUByP+jXVH15pC8R5eZezEfHWjiWU2Szc1
blioW8LQInb4vpGrBhX3RCVza23PlcA5Q0dGJXp36MPlulY7sd4Xs0ZR1kftOy1dlu4JL36H4h8p
Z4cZ674ju47VJ/CU5rKXpOQnu4jupZp5BjO1sBNX0iGBK3zghD4aEjRNdoB3CoQrf0J06qYw3ew2
tOLV0DcfyToJVVSmsLsj0j6N1xQq1ASX72ZcLUPywg/6U16Zwxk8ILppxT0Jek4PfUnfghwwDau1
oPRWtZx2YJDBjpmBPUnTgg18vS6qTQq0R5j4WOsZuTZDUmKRhOJbMbIfLwwc+BDj5Q1meEASl9vB
BwxTZfmLDPCafMbqYJ0skBlpy1F0+CLNsdHu0sYm0SQaMlCaiQKvBNnQhew9tK7ytXfvMlIVgTk9
r+T+6+n7l4nRWLyXYDQBz4PaHsEJ60EBNvC+sCX887VTd4NhBqsnX4zG3x1Qux1weO7Pfie1xvW1
oSR98qYBuA84/89Y+j08oZOhIo4kdx7fU67usflVEHoCF2DDNNmULOL60qcd+74cEHawHSr8cEvo
A9uyZuRbPQCMUOp23qi6Msh+srwDHJ6UKVO6sTWPSrR0RNsbqPcfVG2l3Nl2GOCpM5uZ7+IPn73V
G8fnoiPiEtQHMsE4oIR+xkEEGVGObXRmBPcVxcyJa4MpeMWXK/tVEcDBwjQdUWjFZySx+7KOSRAN
FkbXvCV6SqIz2o0ioa4dqg7sI/5PuBVgYL2RJw/dvjgeAIHbYHbUGUVZd5gk1GYH4RSgYGOncj++
L9LTgxkplk4MdbKIPmFP6RpCinSlx95SEQqQ6guSOEaph/rT5p8WvDvP9luuRHksRtTOY4+5BD/V
DOp+ETZnM8oSd6gutG0/PkNOflk9UKMC7pvdxR0qA98AfDiDE2/3Y58c+ta+r7MQisAQOJqBGgKf
sZ6Xch3np375wy7WXPF2CbaxquYbRpfk7TTE2MZyp8/kSQc4nSCZ/m7DxEgolxJXlqiP/NXnoCJl
vedmAQyCCF5FTsK7n4lJIFqNCKGHhBehHoJy7IZLhruNXa57fkNpN5zWxIA1JZtssR3ByEWTAuFR
nm6+/KmEiLQGO6Cf4x9xcyW/whkBn9PwGZj31ZmiW0uKBjbi0fB1PeJIXeYA8fLcjVzNABfV4UXM
sOo48ztkN9AX3ONbVvREwksnsFXtW4VkZFZBlu13SjL7IEZrSskj5pAkiqSTv4EIxhpyv0iYML0X
zCg5K+foXoYsz06hoFl2LhZmgwX9H18d5DChM29CT4MGVTqx4mp8gxI8WbmIpYM9CkF37GYEsz3N
g8dR7iewDMj0g+nYq9LzpS3aSKmPM0jsB267edyFTBm9vB6I34CxRilSPqIXfqXOt+vzieKiLzID
B2fRjduFezb+02EOkAyBawu6/FEpg9W7rFXhTVwqn6/JBskljSGKHA2Zue3YLiRVXXomNE0woxse
I+hkDuFKXiJp4Ja1BANOXSsHAQx83sOb/E2RJ5pCLodEDNybYH9EfxvU3++Buw8+6YBX69touEcK
cNlCLQWKBJElopcI6qLWZHj69bVXPddnVEeUC6GkjeV88mR1Rxd6un7gUq3Nqrrz/xVkmf2F2j+B
fOtjfo9CZp8HEONWI9xxH3Yij7Fg/DByzi9uTvM0IkFFzt1RiEUwMNVctzlzTO5/iaEXFE8wTsfq
6k/jlQFtoRnYhACvKjbzCpe6bkaP2DMlSVAL63EnI2g24RqbEWI497w3QQJUznuKkXD9iVTAaKcX
5zP0N6VZ9IL42hLuzbBdY8pmiOALBIYjRtX5ENVSvvGN8R2XeT75P0gTgz9uQeaeek+u1ayZsnf2
gv3zYS1JfUxiwFl3dxJgbX0/fWnEW07qkDF3z+0VLspc7efUP9CzZfJYLE1GJv4a9qU2ZDPJKecL
8NHxlNcO/yiR8IAVjQzkJITdEFJ2WHMrBZdBLtkimCICUN3iqkSqX2XrgNrH5Ibm6AlSRLPe46Ky
Gx8p7plZRSASqKIq8AHmmZxaEYtrgd6JtrIHdS4AvGgpP2pvkmhEQOf1Q4qJpwAWGCi+sMM9dGow
pKgqCccKznYRLwjRXnfgGWWAnzZqvlsYpnanOgLWo3YJBY2n/S+hCvGQAM8j3KfJ7w50cOmx186H
QhJVHqsv4PHjT3MaraoM3aT1AbfSamq6N19OJI0zVm98QJWKJ2y14ira6esAzaJnmPEsX1NGOMjg
aRESt/28PqkMQhPX72DAKge6xVJAL8Z6Y/GAqEOUzWieJ0ih7Y6pdWGiI5JJyZ6DvFny9bOBl1KC
tiZTsSI4Xr1bhToLqkhFZfTby74hLC9tu+nPYQoKOBuH78sScjcn6yILQSkKR/lr0CVvzrRHGhjX
9W6VIDjNTDqCydD4Mf5f7WeIW9jV9ncABrM9rSFJGZP3rdmtzEdaJrfMhh7/FxGLhzZr/OrgFREd
ejWWM2z3Eunn6e80+4UClIXqx9R57qUunRVhHzr+NRsxz9H63wrsBbQdYgZjHLHDDJkW5R9l0RZ5
ld4z4rnfF6x8D/A7S3CYMiMT0Rcl/fSTi/vpCh/kbtugIpEWsHnwJYoguuJf8EpVqMQKifv2b8fa
6pWbME1jK7HQB8iKNoTt4kcK3F0k/H2f+w6C90dUA1zKZWuDDrfx0N4QNgdM5sI0Pr6hg0zY7BOJ
lVwhdTdyJUUHwcgcFpJCmrNL2hVM+Ov4bG5Qfe+vK7L8TzjFjyttwEoW9SyZ1l4TDwfBWcK8N7sD
U5EqzRpiruQmwcr77NcYA7lpuJ1a6We0l9lv16oqL5sPXgundxsWZQ9+tEiNCbWtxoDlkdP0cvzx
p8JHpemlrOKC3d170aNCW45vppk78Bg/saJJW00Ltz2kj0jhjWJ5M33xg2ed2iIaRNx6pueQrojO
GUVGfb7Vu82hZKkeN6QZZRlD78C5o3HHKvoBIIYE3gs3VjVymN7MCAP/m8KU9f1taAxnH95jpDRJ
NK1uQtovz4Kn36s9UoPU6gX0ezfX8yXnSy6Q+bjEvuerqJ8BVjr4kH64vHS4FUd6GdAOKlqzK8vQ
G1ZohZZPqALfyORI+6QcLShLSDteCI9fRJNXcN1jXnZ5dyYctCLGX/wxpPpHFsuxjtmlbEt0Vg80
ugD7qtlwlUAnKF1BpSVRUUKklSQrrDpZOhTqjH4tqZ/xVJhE+WEWv5L49z08+jmH7S+7uq1ILnmO
SljYxhNUtULdPQcfVTN0zFBAEBHxuoUrCJZkoqlOQC8isIAcahFHu0YOxb2voVGxPhdc/NE6GsjP
UumrAf86+17jKPIFezuWDiaKckXzzTfsPM/+XrHHyJlTawxmF2Ymg0HJWPDkU2JKfQS/KU1pY+Ph
dVWoAhETB9GflcTJqt9y7V8nRuYVVAIzjkdb6Q9D7WYRI03Rhn6HoO/uXbT4ViKB38vVa9itGH2e
bOSRkZYJatkoLbCN3AzCFwZOIjb4pKgiXOTuIirQ+evXenZ4qkjYHfT1/kV+7ZPIcvGNAurQjJaM
qy4s3ByvfW8XwIIfcgj35aY2yCOPY+cJ/cFdUHaLOo+hD/FE1+lp4cdjXZ/smcjFjxOkjavHPEX1
L4jONIrh+HKXcfaIoMOVfLKF5l4WcU0L96849cbhQAC+JOM9VgyO+tZgL0tHfO8n2/WoIxw+orVm
6D+xGGjfg4FNud59Jw0vYazk7mK7WRyi76aGful4BecYp959zVxBYVM5/woQ4Xo/DFO/o7UOL5KZ
xohQY4k4dHpwbfxYlMP9JdosfW6RrLX1i7auhPvPi4ho1rhfWtDStvBBYw752BCPDKKSd4mgx3Bz
x7VrEaLyWJA7TeBc4pBZb+SVN61oH+q33TxBhc2lrWAZ67yA0Xexi1ivaJdzNPHoo3e0yHauDiT5
vll6dwCidoZBFPWGZOsH0creH5VQj6BVK7/TfjMuAvUEbaaHDSIHNk0h720otHbQU5sxIeNLbxS/
hWEVpBqFr/SlXpwayGKfU+ywpnWOkJRURv0QHGNsdchDGhiFk+OqqL8E/m52ry+KYKvHC07TVTf1
0/m1R2vNf8hxgZlaqW2Q0DEiZLGncAWVn7sulOyeoX++3hvsDMT87HNWkD3kqUWDWDYEz3L5Y+k+
itUxrZxwFNjW4vyvKIbb7++XjxmITnVPFu3Mofcw8UqS21E6kGLoNbbTJCC5E2W6g1lZCUcr9B8U
vvzXbxKzpoDn3Gg88UNpdmj8sfYCz6sLGM5Fczb93x2v2Ut0vNC+pZn1OD2j3fR1KGvgrLQo6Nj7
Tgrsdtnpfq3XZO3LuUFfUPSNiq7yeIBQwFi+4iDhHd5cpH02b1t1HHJAkYojnlP2qp9ofx0LQOIz
TOTgr1J6rcCxzl0SP0Zn+2U0ES3qQyWp1ZmjUWK3tUFL3oPLeL5mwXSk3NsDOlDb0+ynRKQq2OkB
+UFG5aFrM8V7yT0Gjc8nRkHc4z5nlDy6M8532rj3ZinjSfUciSKTKSQUp54iDxohTkcZnSQ27BsM
pQ+r7I2BytrHmHEGgo8IPBW/WrsIYl+I2cXlHsLWCw5hRXlOxiHCQ+XLDCGY7mDoSDclTTTQfeIm
WwT8P2uAgw+1EY1i1NKdZs3OIZUyi0tPcIYFEOyIf5Ea7dpeMt6Al9MByjKVSqq5FMgnmJcEqHlg
2QETbaNodcM9G8qSjJAY274SB9F2jKn9D+MulvZpFGOXWXEZfWM6YZfogrvj9Z+Y1aYWQ4e77qv8
cSK9qX+NIfd3AIUgibrIR+KCdioq3jHq6XsostMc5pkp6mOryGuzyOCMzFvqNewGABqulsuSbfuA
MNa3ScgPjj2J5/UtHY7vUCWFT0S4pwvT80T46ghbOpeopV8OrAWdA97dk0wAd+HBCvNolnEp2mF9
M7IZB8nN2szgXBIlUYOB91zzzZF0l/vV8RuqSOLOWxE8TKqnloSAXJ4zxTIDcXlFd/OyW7tBVQT0
UhhGLide5wJIGit7X+QEUMqVs4AmFGISGk6CPKxnJfXT2wQVf1t1XVLdeM5xvXGw0teqbIvMYbbc
fLEMiOWTdR5m1tmmvpiSj82Q3K7wX1OrkY0vJ5REubUKjmcw0fpviubSz+RiIqOSOCYugXLRXVZm
0mpetDiHoT86fTnCrbCw7Up6qWtNpZGXUaZzHy1FyqaI0Q2KYQaj9o4LwdBMEhiGOBFTdh7XpUo4
5acONoteRiuZB2FXR6+tipQxbovTo7THge/tLKoPM7ymGihKrA2+1FwqdKyZSY2DfIP0KD3kifxD
ZtmutfwLZ/aK8/eQHgYsY5y84Anr
`protect end_protected
