`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kbk9iTSAb/aOpSOho7H3N6ivfZ6qMzB98uiduoncpS6wRafUNEGwPsuNNXkaTQiMvwVTqTjZy9T8
XosdYTuOxg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iwta75MhzULKs3KdshxHW5rHVq7vuoZW7Spf4AB0bfITDyPuXXsqOPbgkVsVVtTQrzLDsL122W7W
N/j/CbNPQisHb0ESU2DSagS9EPBiHpIy7EOhOUR5sePKplyXxUjiyb0zYedZa3+0xv+SnjoQDttN
vBve6mdRQOIAEceX6wY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RDBKU8apkUiOZ7o84VMRvffPUQQKB0a8GENVSKq/b0aEQYMEQ4qKzlYEO2U2mSNGrp5s4LdOby/t
pRqZ6vH4CyNw4Btj8wSKrGXflqYd9Pex+nQpWrIHUlrUubdOtbnvjuqowRL3SnvEg0HCwI/noITn
F+pFI0UQ3zqT3JvxeT+eMB4exyNULiIGNa9+/bl+FITwCruD11rHi+/o8ZRXL8nUlZhPvVXxqWxr
hiESE3bHhGBoctdMFM+ySJAKWsTNcNOJq0kQGAhCG6pjE9R9wAawJVUno0vpo5U0Z4+Em4IZFoym
UPprGjbd93rZqo+WveK9xlWVl5f+CpkrYKP3+w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1GEJBwo/81fTYvgFl+KpUaDW3UWpBvPvi6uK4yPagDQrWkkwmg/w5jl6XzuWpOHqMSZc6InYUN6J
Bwp212cUUfUlrL7tNNSeF3ZEp9850E1GsWm7Zfs1CeRq/myl+OA259w0gWtx7kPDrFyd42rVNi+r
/29jABb5jNsnJaWvWw0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sM16i5P9PM0vp7XkZkMzJGoJf3yakF5idXiWlz6a7SNBeSXk+Ps45khrmVwDHRW++lItHq58sBW0
ZjH3538/aqFSlxlsgR9kX5mhlrHs2MAFHO7wuA6R9khWFDs+F8YbJrGCu9d1awYc5xi2NYbUxYmT
gPwmhIHP/tNWjgk8+QfQQDsFwOoxq9Y60RUGhN5bESOTbG1WltElKfLs0kQIaNumoiMeU1ZJUt/C
bwA4WW+fRhE7jjlF1y61RFMCBeyPmomvwFmFx0wzuVMk3bVYcRaPmCVSWSdjQLuV+ZWRbk1UuwCT
WctyLIoSMBZKNQCBytqAhegDgo5dF9fN1Nt4Zw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
St6zbDRnn5x7A5XQhdmEjfErDnjoqEgOVX/xnwQlArO8HYrEVZG/hUkY5n+j68FAMdbTO3Ly4TMM
WNgqDwvwG19Xi17MJUn7dxkyaHWUih3sWl59Izm0ZVGseROFyRxLLFM9sWpW45M+uWzHSnBcCEHu
SlPsXOxmAhXhx7MQNIZhSchbSjKaIP4BvE5AJSIQNlnXr0/++FOCs8i5AOFDtzuU16qax1p5jKYx
r5Cgjkjou9QNcR/smQ77ALdg69SqjoYCBBQmr90zFZWysTRI6LkXtWOsRNvMbxI7lKEN2790zVs2
cxK0Hb/yIPOTp2FBj4OezpYGTdzEbt4NP74djA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 119648)
`protect data_block
Otj4CrwByxgTD6A3xopEBwO+FLFlpuxcefjlHToKw3VOdAc+RJ+TqMNLC8BcIdbKjoY3u0U6BMSj
3fAWRM+20eoooAMzBaZbUZoeWu4AfiWJAZuNxmSB4TxutwAnUK1BfswwzPV6Qf2/svtcIBYxTpYx
cjiulAStJKPC+2+4W3FUhdGgPqsneIZxS8G3zVHV7IT7Doo8jqtYtiHkcIKF0429hHT9v7YcnhI+
HDN5c+0oMMQHT14Y/w1CBJt2Lo0vT/KWRdWi+cKv4W+FH62aWthHiE466/MlIic6vit918XQmtoJ
lAQagaxNBanG4CgTsiK95QqW7z2mbyEZFPKvQmVNETuKtAXhhuC03JjklK5LTHcTNuTSSrbGBpAh
SVFO+mpalf4VYWhbdtn5So7h0C92cqvbH2RYhz7ub5Drcxb6AnZMA6zkTbt1L/ud/4CsbVBSJ5HH
Lj7n7uQQoxReS2TB5OqzjirWtJ39tcZ1hcYAk8KhLPRBWuV/KQrKbA6b0i25A02kh8ll8ddrirUw
35JIz4KUkaNcI29bfmljC0ELFVil6XlD9i+MN1oTdeAAJ9U/TgpUAdtiqiXM+4VGgaO8/kSF7bC5
q9CiNGIwp7K0GfeQpSycb2Hwva0/y1eQzY9rsbclEB7cldauP/fAoKjoDif+iiyHVyV8d8YFxsC5
rshP8HBsO7XIb606rbu0AQsEEuzg+buDqcUCVPa+asXhbuldxZNBoBqFOB3V6y9c1jZ3gxKWrK6p
fbiyvV1feC5kHPXDWNNPqTDrpihKKrl4bonUSarmlmqy73kBbXXkDGW1EMCRqLohDzMh49VgsZtD
NCWofKCYUQlwSWz3upfyRad140vNQiex4t4r991MIWCXvuIN4Qyw51Rv9X5qsqLVVoO3KcUZH/fx
DugdA/SApRdyb+RrRQ8Rgpup6vaOINu3C+GJp//Pi9cDaPiyuRknfLtRNBLF2d0i/ON0heKQm644
p4kIzu48q19Sy4oCv6g8G/UbmTHNuM/AJdU9A06Rh5/3gXOF6vbk9Zd6/JvaB4APAeh/sB6aKZBD
JQ0C6LkluknbuxwZRYX6AhwvBYayUKREW8nmZyDN2lBIU9UrSCJgHbcy5y1hqiDwDS+6gJZ1mcw7
6JGAFnEM1dTAx++kQBKfqBfxEl1OqNruyI2XscQiZIXbfAy6EnxnPWcbTyZwg16Ev8TQqtsFtUNJ
fBSGy2oWpvf3NylVVZyut7fyNpFGE2PMEZ0tYHm/gb+s2WSGhGAlU4ckq4my3GSxd5gk34Q2mgFx
80Gl8W8UlJuPKGFluygCnUYpJn1B2GXCtKaj8WWJ1zaWD04TK/uRnE+d7oVKxlKxaLktAgKni7k+
WsATU7y98AeHZIuNKj7XIHt4erqzMKPkR9IeoPnxi9ZjxuBW8OGrFV1CdUYG11JLBYLJ95PTdxKo
JEt990ZpXm6MHnL7btgR14jjOfsmgBKPudyjkpjZKhRAikVPOzVkuuE0giKhL4sD+5OFtibRIA/9
OEfHcHwb81yJ+crG+8yI60BjvHSb5aDQGxA1kVsDhuL4UJrPKGiHqiYkB5aV2mkFPqxW5HpaIrzE
SyE5wvzkk3TM98vBssu8AMj1RtImx59SyIISU4GAybSTo57wbomRIBtAYXgbwTkEbxLsDu/PilbP
yzc1NQ/0Q3hj+Wax/I8z+DER+dVkIcXSY1Sa+kDYIV3+XvtumsL+ZrQuvhOPSZu20lx2IskQfk6r
5olZq0xFEpK2mzmDnhPaMu2JS/wPnbDeiP+S370M+xBJ3pytolVeKuwYDDxmfTXq/gLjNaekFt8K
1Rgu55KmTDPwQRVXCKV7jfmv7HCOtAkS0YHFX8R7KVG7aGkcP698JVZhLd/eUEDLDqDsUnUswpAp
luBMYwBCNG55yy+mkiX9g2btqK59dHzxJd2F+p/AKT1J+zLGWVGwku6/aBoWmFUIPYpGV8EYGL9w
X97T4upJpLwOialKMEWlkshqFZM9IGDGHoNE1/49AymQwyqW1y69XqFU+GTrIPZ7Cx4APSPtECaO
qam4peX6vk/rVi8XQ/KFCDXc0ftkubZw0ieCFsstiP9RtGiISi8v8pUeopms9A6roDY9tJRCaYeJ
bYzwQquOQLioaGDHaWI/OmSQ1o/c+0nUXk3W9A8ktby8D4/QysQgHEGOVQnphfWd9KDlH4mBNDn/
t5lI75fbk5mH78YKOg1FhnOIGdtq7YzPY7+l7iOpz7Xwv//LFOuPypoOb5BivK2uFDtk4X30LsMv
EXIX0uaay7NBGtQNfQApYn5CWwwavhnK3QLAKYLQJ9CYAbTjldHK53cHqQRmwpEXwSN/uofrF2Nn
JFeSbOH/dcqNuh1IkXHtBFQhkrsrivgSQLl7jwd6Ea89YBwfST1La6QDUsd+9hFSbTyKX6FquNQ/
7CS+0Z6/GIS3MAzZKdahVUVaQ570QfDp1ASjfzzqS4/GajmdTOI/yMJO4pvLqTX6MPvl0CxpMsyG
T8eFznnwTldSJGDVGGhBenIQVRZp4VB58ulN7DTTRAdf3oEKMiXhkBxv5x1n6w48V5dpQyKk0v4Z
CJ9Rr70HTWpEv4OiCh9HWyyjB/4qW0lZazwTf3/EQwYXO9legqLWNjIGQ2tNBHFeJqoVVzbSx2/p
Y2taIjt44gye7fM65kSGZA4e4C89cjyG27Ji/rYGiMvlneaL38aarDbHALqJ5X0XLFcUSdHFMfaT
wBAyk0dferyqheTHsvDnkkfEv7cFGgyka9CTv6p3UFxQWAiLIVlm34pXhwsxw3gNtH2qNRtWSc+w
vAPDvJpESxSzFi5kxGfcLNjEUkt0PG6mfTs9KeiaaTp6YfmKGmEy8n0tj66l5PYWYVVgtFppeBdP
eGWbGnIX1z4EtqSSp5Zy2AeiMfZ6JBZlgEGSFJkV/rEADKJvHBZDiCHy5Q55n1jgK16boseZhnXu
U+EXrFdO4GExo9/iJQ5gXZy2QGv7S0azaBtV0QkB0zqBkVs0UB2gWG7IrdfyhMDWn+l+uW23NxQt
SWA9P0dO5zWhvP2ldyKOY+rMrkOMnyj5UXv6GvTYeNTuBTTXfjejbsmHt5h6eHTFUy0KwalTbSnC
toG6mvDjW4eXLULVGyCL+HfQoxbtI/57fTHF3+NvTazCE6rs0L2N870Dk4LRErPcf866XmRy+5jZ
Rv7Gf4WP8QG39jxNa3hjpen4ixeKIH45KuseCTZvHupkwae0dMID8I0nJTzy2FKWKGSMczzVD0BZ
wDSoQ8KxKdlLdn3qzmuSPU90eu6xW0Hsb48lhQ/djy/kHnFxtsBWbAQwOEIO4eeeoVF7h9DMVwbr
AsfObTUe0b3SFnCffWA2e2OI1SV0gGZStA7dDVnRDfE8u2KbfeFM8T2NxF5pHZkzo7UXrtJocGrA
9FoAJePI4pYv684DdnRCMcJ4vQiMLq/KvPISB+8GeMzDz/G4vnsv0ED1rga50ejV+TFFOttkO9k5
jypmNxBlicrmdA2SjXuSHFffAv0/gJeYa86o6j6/UII6hUGW2fEs6bWMbiv3wMfqaFqKKuI+v2oE
m5orM0a0cl51/9ncJUy6qIJpBCI8ZK5p7JFVNQDzAB9pMYXXB6Jvi6ZTPWf4erkBcOxI1efvUQEg
ll1s7FPlZACRjMW6wC5xvADRwDuHhbtTJKDX+Rk2eSJxoMkjUSMIx0wN7Y7NRmtI7TmdK+Gc3wJC
dV2YiWgQWmUKqJwfN4xXo3zGXPZLbLxkcZMDKGpnYwt1R2Ua1VgZuQepTgDbLqofHI2qu9dgweuE
mw/3Fbw/WTNHf8i0/2neMW5ml0pxah7OOEc+TzETstMsfPC6G1FPH5zYRr20RO1pHgA8qLMOi7qP
rFC73+W5EOUGYt7aSlr0jZ/WIEzQ4PTM3Id6SqM9osetcHqzx98C9VmBTUqGRuNGzELhL1qdmqgA
wDEWRGKX/kH5ADJ4mS+AxhH5c1wQSQdJGdtvWpYcJUJnj2KgLgocG4jJttJPy0n4uZcndCiokyER
TfxRfl+YDV4dLdZYQeU4WPwJyAMmV+RnvdD3X0rinvhi259mzXth2z0wuoNO/xY5qx6GcmGnnayG
ZY/ulqKE40+m4Ha+pG1QSDZqXpsuoORNkaVuqTh2zVcFggDH2L6CPaeRtp0wsEYYvk4ylWTpgJka
UGaha1BV789Q6+mT7fe6GscunlDxt+z10Zwiyv978JhWD474GTkhlQ88rW4c5RjWTCVE2MhV4tMX
OPYfVv1rU+cP7AcnBqzJUl8+/6BKzBESApkUIvMv4XVhKiiA3AfeV506fkfOr3Bu3jvSYe+anKyJ
gXtqWQ4VQmWt98y6ZLv/Q3Qmiaw0daMaQSH4i/Nm2RbwXm68FJ8eYHCkHVmE3BSVMc1UZgER3FBM
q9jMxHe6fb7Eac/GPnHdi0CdADxUOp5/ZzkBerVpuuHP28ca12jkdiXmfTyQ5s1YjB8jIm3Vbe74
g/e4W3ZwfjfNdKAiVj70GjL2dI1SxniKamz4K5YwQ8Hlx/CWfXqM4DTNViKOTHUF0cxZeFLcpEKR
q7LX2Sf1ePyhYxwJ+d+DLcJKdHpyxQWZjb08cBOij5dNzawLH+n6iyKaAKUw86y4xkHaA1LL/js1
k8jhWba8Qzqb3xK7oz1x5t+Sb4BIo/89UWeqKK5f6CoaKY/Zq7HQC6GLPSMozvRO+brCholyITm5
eQTxO+RJHJxmNdvd9dta5KsBWzOh4B9iUxYfQAMNrqdgwT1tOik4u/d9nDveFg0sqDFZfEoB78tj
hVEJrh6xgrKQJPWzp40glnZ6/wGPHho4j34G2ibrFtnVB0HCO0MKFJWH4fsMJMOVjg8YgJ5rdDNT
Y6EJiZxNjn3xsQM/8g2hRMTj1PDlQ9hk4rB/nHGSsTkr/DvoamCMcggEzdpfvwXsTfZHc76qHi/d
LNKfYviNifocsg54UjY5wONVMRtMC11Kg94f6pyPC+2oLuxwU2KrAe/1AGXCuJ1w/qmV5T/QsXCw
zU79JwbcRGtbiFSyMHMpFvq9N/dVdBuMHMigPRzfes9Y68pMeAoWspCPW13z3vZlqbrHqh0DIca1
4IU/XiBtxj6i5fvNbCl0rQxdrhtWYQrIOe5w+y5XJqYS8eSBVhsxIJEOraUqD/gjpXl8IyuXfuop
PoUHAeUfujR3Lky1Jlv15IryGGavy8P9mUvTyNCtlVLZKo7aR/Bveh8i6szi7CmhP7V0KoE+usaD
E1GVmjESHlbiXkmlSUKp686YFS71MtLPXPydLAnOSi+MaHuQTB/WTWyTIS8OxlSRrCGWvvZuTJxP
YRjc4YkUwRnKeyeJSqjWBHzHOytqQGvnDL6fs9rfKHe/O0TyvOx8d7kPPxnhLCS3npEdbhHaBAJx
8fvU0NOTAlpLmoPiVGVdy97JANAierbTj/GQHCwVHwCIYiJi74OOBH/ZZBVS16nkGu45YAYhDGvg
6icXO2yF/fR5SomWjCEbZYhwxD7GFmAw5wfYvP1Y5uHWqlME0EdZiEfe+dH+9pi9PbR1HD2FrXp2
N28ih/zmf/rmIXffGiHjnD6+UKf0zz4sEBwotEsQr+NRMbPWj1P9++vHiCCAH/dTxMowZNTrEYKA
vWGCTDBn+nkI7wkjamRYR6uCUdlfg4oRdeAHwpiQVdyCzoXH9c8b0HMMae6mq8pAVbt74zW8dyfZ
ec3iAwlEPdsUijxCzAb2n6fhF5EUVAkqOQMMmI+kEDFYokqLwGrhjk/w1YHkKf5NbjxdBcI9uG7L
Yfdtkbr/nO8L2mND/zAn8L+VgKlS/C8G4mEnM8Rx8ttU00ue+kDuL5F6gl17rWxkuZUzmp8jx/tw
jwMBiwKscBPOr2x2J2IFBCvUp6sV5jcFI1ERrgiYI6Atdsf4TVMtnuUh2EdjFCUULZBXM7N6rY+i
jrJXMe7/ldU7fG+cDkple0ZC/0ShuEUDTA0tfY+EVk1IxsWbWkHbJRCXHOFhTP4kQnKE1RKwpN3t
w5seGamoO/W8p02+ll5bzeEwRrSYfy4da9H99eVAMCrFxTvLyIZdtHarbinpQFgdOy2c1pLfxUau
hfFn7XgUCCbha8owi2074mlJ+d+yI6mtCtIEGUE/D1QMnXiQ/CMtCZ0ftXMJWzQ48irnE1lyLMee
nFuonI6oGA+CSrtPTKjhG3EOFV6/HgrTc589wfcgFSGmg6wLN1Ssu0IDB+STrHGVUlOpMSU5ObEG
oB/PH/0CkwdEoY45Y+kxBM0dtdpqtUxON1kLckOR6a0V78LknHOjMsJ822Y/qJvfOzvRzkoEJvld
vhlh8uZ7ek3QtcgudCPAoA4SKkLzRBfD3yHJOWLpgF2cxkCiYEuclV65ACJ4c1Nc8i6JfWy8o0Ue
o7VVmAHmSqVKpZ/N4/PAUch4JNk9iNJ6C2ws/w6HKM9GlK+UpeUumg/zvStyiP9i6+e/v+4rm1O3
0xa02bxlKHlj+4ptmW9fO0I1VU55GvOkSot+LBVSKM6HGdihoG/W8/pdziF7KMaZ8P3ZkOCDrzDJ
8pPcBB1z3mVwDefbFw5qzMif/5jJdp0pMpxf+sBJ/Zck+K3owLZF1OY2qqInY9K927KI+QbRG8lL
aLLk/PJfHEiofYjKWDSrYE4pYq5HCEbHONeGizYx0rbQL/mKYf5gScP7u9EfEuww2XYaYbvFoci7
bvmLJk30r9o1fsyCz6LK/nVsejtd2FVcE8O2Whwi1RqU4oNXWvE6JQ2rz05VjsUSsy/W7aFwceOF
PUoQQlwcMVmfuOVh9iWDxB4vnnKw+kFWJcthwhTsjFCZVpQY9HfAVL8P680XH1XehkklzURHLgEn
KSxrMGHNz0gy659bv39F3pAD4+m/NZVjSnH/h1OoRrr7imqJ4jxfyTP0SZxpyrERKOFADBb1fc8Q
jh9uqLBL4JwbM2lkNgROiloq6z3VrgvciA1kj9mCLnpiCEvSkuw/GOtQvA2hiU0DarkOOWuOOy6b
uTpmD+8azmBDvzXXPR+tq7E5oBGThL00arj1/pp1ooXaSSjLLKEnq3BLa12dXg8TA+Vo9cQBOsIL
2BiX8TU4io+vGVMhVvLsrg/IJjZLyxrfoFAITT4028au6b/c5tiQ18WWTU7ZPn4KYcMDVkjdA2/2
Zl+Lm8onMB6W2G0d1Di7TP3mzhpXcLcIm0er68C9KI/zu1l9bw/ZWFPeJv4XWubJgcyIhgj0eIDT
5xGgguVJRHPqbOFsS19HemMWUmyr6EBfrUGLNxL8NudJHKQ6+geeMw9YiPsDLcUjXrTw5jqhh2RP
h1arDcHOtKTkcvjyg9KtW2KrlTU/lo7/Kduxepql6ERO4CqDnxw2w9IoWfJze6VW+wcPiSzWZDpW
/lcA8O9FVWkjrDMTA7rvMUqYAT6nP801GfzSPgUCHXVqS1UbL8YH2/rYVvj1uyLeKn8phUDBKSTb
D3Vqs6tmzj5ojIcoDYGFn9MlVM0hdY53nUrrsDgEGVl6H2QZ6nZzK+QoEvPEejBZrA4j3IpgAMCs
IE3/C7jM6YET2GsOl8JxCGQ8TAIrMlIG1iiszYqgDkjOUPKjVyKkEbMLKiKOP8aRns0QEPepKoKx
vaznYAzs24vj8OjE9gAmSaPp1vwqn8TGjWftkZlClAKmGrEMAS/aGams94QIpx4eZuI/nNqeo3W+
ctBmwz6/8iojqkyhxxXNa2rQHaRGlHbKpr8Ny+KQK4/cFjQL5bkPOXM3RT90gvRRNCHQ8l657vPL
4lS2Y3zKD4tXVcP/DBBCjfdjJsWE0sXUjijQAX5NNvqMk4NzYjW3aEDyvxnHF8gBBEi6spb4Q695
meK+Lv8CnLiDw/5InKfxmdS94cpXCShf0F/YqBs2rgLZwXMEB/uiUgV6DE7csR4qBTh+1gpEab0L
n6pPTDoItK+bfTLrxcgf/U152WS3qice+/fhVU+utZCCcNJNqHWi0er2vqT1lgarHU9MSnCB0JHk
Zeid7eZ+OvSz79PHTlc6pqc3pzddv6d3RhfA/EBd9WcsBRMufw7SjfpEpU640Hk1g1gg+Zm5qLX6
abcyGIYNaqtVx2K8IRYb26QhPNXuSRTCr7SyXKQhJNGfLUFv9LK0Lc63sWTEk2mUugMgrcr52Khx
6Ci6bgOBbljaU38G0PyzFvQuBq4+0B2IRLJKO2ALT9TMQQjjkXBzdlAhXtAlA/v3UJSQSPxw48cp
H3ZTUkDNkQQyAkvHib677iZN77RhKx3vtOrKcrAvX9GueiKesbApyitOeYpWFvK1sShGNGjQdfgN
b7C+/J37SG+L49BPYe+7zy6fT7uUI49b/V3sEOPgJ7jITH7vaboFEgSbwktK7g3ydAfVO5+KP/HE
pd0SgEBn7Ww75fiPPsKBW485Lh2TTbT5SYbnrWpJfgli5NENQbZjA5cDl9Pq/iqzhJi3168HAMLZ
bbwLoUmdvf7N7PIjbxPhkH7MSprRyUFPOqKoX9uiX4Rk1r99fYjT/inD3mOTkqfJ3O5N8uIy3wmJ
VTCvhs5nOY6mSfmCVSuyAh09Talw53mNmQfHKlAuW6f+2p/2iPuUJjL+dN/pSCQtFcBylqK7ovqE
EEwE++A+0nbn6CPMe9REqmY5SgmalD14RBzaBbN9a72qT6opWwejsAnU9KbMfO+EL7mTd518RP2n
YQI4b/mvHx164B3sftXx1yt26xwVIgrQsKwkk/UKdqjfi9J4e0FeQ8223U+RTTaSBHUDkaUDyV+S
90onGBE6LoBvRYhOVIQM4aXPoSePaTdLqapPAZnWsstSpp9Q7iKmhoKnWpPORHaB+45pRpb/HVdl
k+Su4WSv6NZz7eb32LhiFxOKDXZFxF9lKgkRzgi/rVaU903pkJMxllHNcnrHtDrw6UBJ6Sl9kJoT
KL0nbgt07xemRB2TuwA5vgZwIilyxjpQRTwSIssPMTZY8WesBtHpTbZuEBQJlhkPX0dUd0RcZSM3
E+dWEcri9ZImfKDSjwuzC2QyUJFV0lDwu/NHWdWr37j+BemG2NTqaXLoMpPf0emlmvEjz/U+r+jA
09uYblXVtiWQzR6glz3JR/kzmLtrNBKmgUPkjfd4zCPnnseZPHAI0YynJMVHb2EQsi6pAdJm701y
6ypWh7l3ubTQFqynV/CnInx3H2m8lWws53HKoLPYJFpK5HD4sfHFs2tongopOOZ6n3YT148E/h6p
F60Fh+cnYUWTOIn4l0pq5tSWwVIPbcVSVj0twsJD17oikYYkQ0sXkwzx7Ll13ci2e8PlsMeRJ0+R
2gyqqjUiAjZP4MyPAlOylNX22io4DSXO2zHv97pX1EzPuXlxBU6g6IMPgaJ15Jpuf6UZA0+RaCpW
VHuv5tGdktH00aSizMMtULSBDA/68JE+wZnVfa7lqK9CBDrpC5ATM//CJOlmofxEYpEefCh5weYa
LTgKI3xuayYrMIKjwQA9OPe/9c5plK6D844HUu5GKlNNubn5hGJ8TDLyQARREBKFn/KU0t8tW1JX
6AhcQxulPVkodecLpPK/dbobBgL3345C60BZGZ3mHOEtNrAVk5qxMG1IHgw1R1BxpO3cN7ObmDlQ
VshFa6gcWb8tWvS1A3VXkjHFhW/m1bterfKjoqsA5Opc7usMZEhBe0qnC0jUKbHrlFqnCW6MuQCe
Z9ZTX4pdALl/VIqaUa9hyz3aw+nmho1H0y3Keb8RQCSSv0l2yUXVw+SHx0pCvmaVbNRS0mGm3Z43
XXguQiDVoUkd3o+qYruGNlc1V6EFTKZGZAZAyZdKogGuukWiVfjoVeW8JyE1kzaduNDA9jTi0DOx
V2JaEmdTDJRgTUCDO0uUDxNNXwF5i1g2RSpB+ncZjT7dDi+AUFNKTqhPt0xrvbU+tHvTIuglk9vl
5PwcVl4wbYuBAl1Ch42gDI/zLNPnVZi6187nbbJS/rZhb3AywPpwpCL8TRp5txHO8nSUNHKrfQoN
HvpcJepTyB9Dk+L+KdverYuYQtK+1Lfke/F+0lFkIl65r2/eUZfAnCV/HsoSL7YX2VDm61jIsNYQ
gKVCixzZI+2ZRSTtnttjklN3EW79D9skF5Dw79a/Q5d9OSNxZt7Gx+PKiJN9EDljOKruaBuPuVGo
E0F30XpFSxBd4rFTgj8L0T8HQhrzf5qyUstRFH1J57HuGpRN8xploqa2dok27rfCNzgNHdEWhBYa
T0OsOvlkk7Ji+wjCbhMH4zwGzo1f1ka7XD91TY2VUXXxZ3nfXVzVE4hEQwTqYGIkcids1bKUPPZd
BeEkw0HcP9F3XZDMFxZPWS5z14EUva6X4qyNRoNL5hdWto4IvTFKyHp8bRoVKb/Q28F7ZTkaXdF6
evMsjKTEJu+5mRnetofsThlIgJIDZQTQtEcwPxj8NBzernQ1Y75qkTS1mDMVv6Exi3/r0TBk++R2
mfEm4GFrfZmaXBirWooXr4SZRK5HukSpWO+lO8ENc0Yf17ozLf86aoQP2o6jKdlxq+75yHKMMcs2
BKwcywX30oI5TWyVSNYRGzSVr0mV89u3avaWrUY2tl21kpjipynmtFrY61l8njvaTGjYZ61j8E2x
c+AI0uI65QttABv71ild1w3O8b5PNGst9NB2XrbixodqC79QYhKMsJcK6qHeg11dKZ2qv1Fwfn6W
zOwCTWar6GjPovOjNuL7377jyH0FRpC3Eb66i8t0+/P4tiKSKJp9ff2Xnwu/7ZzdrTyGiJp4EUbX
siTkxU0WpbCmvfuqNjDc9ocqHmpkWwUaGzkBY8ZaHSBleVV0v2GW1/1K/7JhxRWcnoAzxkLhzgPv
mhxxKoROBjfYOTE7WzJigA+ZCoR7s3UM+K5sbUH8LGn8Z4d+l3CQIrLPBsKlVfbI2oGioSyO227X
Se/2XneWbOXJR0kZf03cHjQ6qC5TBqwRIlTWf5jVX9bT48KQWEHAH7HjHKHcCweOkCHfAYQNXFr8
QVGcryhWdvIcRrA/aBrBE4LR1IK+u+fzaFdvngNnkVPgbp8BRriWxz6/KKpx9GguiIV0WxmjFoQs
7iF0AVXgfEz5sSUzhkbwgQWQsjLpI2hyUeT8hC0acU9yBe+VcU6tXByZ98p4bUS7QHwXqvKylaIA
dU9R1z5/CdZ++JgQyU29CsNo6kXiDyuJSunGwCV+SO7hcthROpzZ6CEVPr4Ms0znFxCJ8BhP/tVL
4QN+b/+DPwvjWvtf7KFx5fGdEsefVrSRDpjAucOyxR5XomogARMhRqw3N+F8HMKA0DdrrqGDNPBU
LJmEFv7mWuJbCSUHPGM/rQFfRegB/CDAz9ec3LLUCwXxRuojLpZmUj+jmw1697E9HKEqeMvs6dhI
XT/JK4xxQNZbzYd+MZRpMUGBJSu30A9K0olWNXk/7R2OD06qtzVsarannJjiDzcCfN/hAtVEhsdp
2WGgDkpeN3Ag10e+iPdFwlIEgF1Z/i0DIdx0fVVLneejfZRlMFEAfAzE+Hg9WRQJdWeluj9z4kkS
tKCf9EheA+w7UgKqxyMTdtiivqD8j+LlNoTHKvYB6TijjAvSbT0vE6j+YWTV5qlGDgNOrjzwsF8s
0ay7rQwlXmRA4X6hMTx0sc5eh7Ls8i1K4qVIQ8YHSXc4NKSalz+j3M8IrTIZKYkHaHxooXK0u0nk
/KiZcGBQHSG93G7Ju9I5Ri2WCKAiJQSSwVOaNW4xjTD49yPbFUcYhLw1uo0P1kBB0HN1qakYoWh9
suOQXzPSBuD3TEM3/od5N7Eb/QHX0eS7TrqCHjRBxaP/H0a99qrhP805ut+Dob0UIb2Brk1kQGf8
cij1CEmxjRy73+A47Fx3L9Zgc1IFhmjTyAMDe78z6w7p/u33b4/uwKO9EftuWFL7Z9bQNa7o1POQ
DxiUy9Nr91Qh8DhrtD0aZeomUK7uXg3ynGk+y/P5Ad7w6JqeLxcP09ZDtAatwhqEml6thfqOh7NA
QNZUaKmjFnWwgSX7DuPXBLnTHL2dQPGIppEfIHfbQDn74y29LtmQMkAaJMlWWAq7gGvMdnuVWRce
r4DuuRSiIrWh6c8WCFzvweOlY1ppQbgJD5Tl8E6LWNBzK722PoH5t9iqfgMcod186D9yK/KStCpj
PG27gcYQQTC07FmdUwXvW+OhARvgNIjcAvXiCGnPQn36DsPXF8Wykd3e5AfLMNZe+QPUgK09oy/E
HHEbw7W9CGIjljq2UtQFObnqguUh5ZYmrNcv8FN5tFaBY28iouKJaGi54RK+QqzfiN3FCEmVnJts
F2IO8pJRx3dcxh8iawI76B88LSiQUNfMflr/dBy33hespI+60P8B+alHzajRthAy6bRK7eP6Af/n
RIkVjVO9cMQPVH11XSTnm1V1O2+3QQC1QjSvbgg8HrDwZ73nQtQO+g3TBJBKeLN5t34f9E4eIjtw
4E4OuADCI2b3gpNR6tBbdNPqx4FhkxR4Oe+Lq5PK9OH4WW7HvXLVyRzIfTauFzDHdQGC7IVWfEY7
GkNzU7zVAyJWGBh7viHe9RS17X9MLY2dbGq25Kqkur3iDdugHoc3nvF8YaVLoBs6fXppMIyTPjyB
/l+sXC9bsvzuEfNOyOUgFPWOUg32+XVMVNtSBcmyYLCGd3kp1iT7wJp1nGFZyWXRxET7q82Oo4/o
iTX54kshALymiqkV7z1VEtHpiTI/ICxTmZxVbSOLrIjF3kJbADDhm2PCDt+Acf7fVyYsiuqvmE9Z
8RXtVvuFzXZ/61kr9K03LQoPPHDWYHuXzR99dheuI2Rww1eM2EJscHHYhwpi1HzykArmpP6Rs26u
WPm/AK45US7TrTOQDaVIufXpwI50hgy9Ow1uZRYvmBNtaUVxAMOwLnro/vhaeV2nWfEqRaTaKkEO
9V/yqXNVf2anKCUs8GgjDwKMGe9jAqHXSCwcT9Ap5nUlHpq5TPvzQv5fOe+HUIBSFCCUSj3z3uX3
F93M3XnGXqlziQPJ2CHHSc83sstovahsfFiGWhxTOener+cfPhFbhQ15E6dN1809IBbPtB5eHLv1
VkbpLFqrPMzuRLeOmKUkUrMHYv0gvIMBVNymCEUrtGXLZO45SszCjwcsyaFAZpZ4UeFmpEVf0pUi
gWm3uYUjasyz1gd8k9QqmJ/FCuGuQFAWToDZgCJZ36iBRC9Rfif54sDa/cFj3LNRrPcyGEgHJJnG
87Ole/X0dccUfodFPzdDK0/YUsw2TawjQvn/SdSJi+WX50RRXE8sMzqlbzN+MgP3Vs4wsElVwr1z
bqC99hVDalATyYLKvLOGKOxagBfGCyfdBq1IPJM0W8H2W3DTsAkizVkj1ORMsNQRcidY1Y6LV669
a/F+HB2ox3g2lz8EAa3MzTi5X4QOYEiVJpmRDgzGj0wTbkUEoqbKA8LsjHXk6xRyKAoVk8QNOMo+
FA728m4UZIuIc6soxWcMf5cTPxGowt0lGEuzaKjygrvSNowD/n15OWf9zX4mjMoZlww84iVbW7KA
iUKM8cSe4HlSLTXS3CxyiECOvyraU9lDMwuSJ6TxDQHeIltEjaFROJt1C5H53AKv90dSvsUt0FY6
21LysNXa7hZZ51j3jvT1yitrLikLB5Zn8m1AZTOhVw5Q6NP7JZUn76VyCM3vqY3Klq17p4bGwmiH
wOxdLuNBLsy+Kc4j55QBuL4qKgSYjc8fNs37n0ujgAQdz7VYRX/EbtAWf2EeKpEoJ5qiKV/5jSQO
1cU/79IO3agzrePGqen7ELUiqqVpcE5scipi0lNMbx4zlHzvO29Sx5IcYLuOGZ6/HBvzZGmrtJwK
fOyzYZdzh3VfGQnz9KqIu7qWVkhX3ImCXTit6kfOe62eCXAPQIwwqNc3LG8V5fv0fFaTo+aOJHQg
Wuh4wh9aDxWAZMpg3o70p9BqzX40QN5OUrspDoGcL1o2Jfs/Z19dh53djukwAIkFKvXi75mY4iBz
1kgewuNHZ3NyHhtaqmxUj78ozCvPrGersjJXfn5PE4aRmUd79Y64vY1OEHdGzOZYtJkgMTdzsrB8
6QwD9zq3mQdZX/ozutE+ZYHDecGHbI53SwBFKWhM9FOVBbK3DSOl6Gm2eOUhRx52xOMnogxaUdnK
ltywLEk87YmFAc81RVIZrNPFWQQiul9OaN0rlyxHLi1kRha2qUqHceh67f6pvzlZ/fqlszJVl7oQ
DmW7N8fy27+JjwRp3QBi05w18baeLNw+9SDgjQXBmqwT3i4jArKzuwiMyZt4k/d8HnpB548ISBZ8
ga3SWsGC/O7zLxPmDxL+ZaxisOClJfZaP35dfan/3KZpMUU3ruPWnNL7MJarc5m32PXf0X4dfsJS
R9tnkfWHNFi34XdLOeFu1KPn6utBQglRN3Rw4RJinvWgIzVCa+qIZFvlK1qWlDlLzikK0d2C7Vbt
ejbeZHx+CkJRresQvT2Zl8q16omfUI4yAendpTt1t2p2YZ/VhXE6NC4xzdYwTarPiTBtbkWwpGZn
yBb+ssaOs8jEv2vgbgqTAB4DiFe3mc7ncS9VnkCu7An10ewb6EpSvLyXTPJrHP8HqONMzsnTxx2V
MR99AlH7B16q0kAsuj35zbjviA2LVGDxq1vmkDQWKMWhgF0xePhU2N6vmQu5vVtUxtZ/oQEG+vhN
2WI21gfKmQdB1JuKdYxT1xsYxZVlERlK3aXhfD6Bz0nGnFAKRkUPtZ4m7V9pnLqkylnwir0/ItKu
btingJRzCMu7IME5UL8J4lj5MfdzH9W4OcX6TznM607bu1mzFtdoComIclnTRDmxTtxVvrfPbWCK
hTzU3/Ks8OgC1UseaAyBGu1ezBbuMYVTdov2VyFygIwDbc9XoN4TTKT4Jmealu3N5/L3yO4RLy4s
5f0PoRRoW7IPkOPftuzeBHa3XTpMMWVMQd/+MePCWWdGOJMDlwH5o52NWoy3tVabkRovcgL7WMFa
MEc7j0oeKMGufWt5Yji/ZlOp+kBT6t03BbonelwVKzz+kzzfYWU4AyMvLcmg4ZukV0Edv22R2UQu
XvXkQI7oFeria/HVpI26qSpzQgRQdO/8ed/lhyqFugjirfMPLIeP5PdmECFPbQ1UTuMxRP/n4GD2
0RCQb1crKYlXG9/Oyk+fREnWaAYT8K5+AoXK3erqySbms/W76OSUbN89Bq5UcxgF6btPnXwrOPao
rZb2Y0VEc5Pa/y/NzWeRDyHhUaUY+e6+NJGmcFuhL82PQ3aZJG6AhjgCgrLvKHlKnCXv+Kmgec8y
hUVgWAEt66YricsJfITC1YAd6pu2iQtHukkMow6hyWjzNfC34Jx0eS9hyy1yFiPhEAzX6XCgXE1C
zpOxKi9Fpt1Ld+a6UAqMjTLCx5EkPhmdE21PqB5scVJYR5yfJPxiMZVd9QdhFDmAdf7prmzG40wp
eYfe9UtJnlLW/28FAYXizv96DpFJpcbTgTLgIm3ZzjhFMelsjH3MAkqG3aU0AQgssgHJaJ6y7Apc
SK2fpIpRi1sB3Ud6uqaDI18xOPVnfy9RkCJsi1UUWzMi6bmdSR+yJzrD8d8YraJE6rL+89VeUu/s
dZz0iMtJEexYvZHc605mOmaGJ62Ibu9GbqCXXDmyYpoKOgzqDp8Qk0aPIyGJQQ4Hayb3/ffUhehh
zItoeot/S5lejRsWmfwPm2Fr/9LIfd73UoJFVrdJ9qJS6eqk+20HCg2fcyo6zyhd6QWFfw+ilPI2
AmIG3gw/ImzBjU6OyUJiPGigg8vuU6Fdt9+yJ2evl7KYpLAD2Z+Wqekx2Ev+VPSxzm4fqm8ArrVx
ZK63RbmVLQWZbh/hs4hVPVbNqWs3U0nCbAKoh0m0aUGBniibB2lbReb9JzKY8pYa7mTMvXeFR2N3
c3EwOvha7tFUs/xTc1W0iSXXkgOxk23F9wwY+pkbmcq9cvdzaUEs/yp5qU/sjwPoEeHedCP0leb5
zvy+b9yMm1VYqxa4gAWs5jbValolEERbXa8X2JbMRg2WNViIhQl9UBL9nYcOEMj756/4D/rv8h2A
vM2fT+7jlGuQoStqnOmen2tWzEWFok9v3hXEudbw+sKNCGOTi1omuGuoOCjsNDgbcMmrRXjrUIFV
pO06mboFr2XBJKhSNEkg0VLDt/gsn/6k+zJMFo15SL5qj/avV7qboG5SwVfpQslEXwFShgU4yB54
3ybOhmHDTZjZldF6VGEgEwm0FIeI2D5ev0TvNSZDVM3eu2+2VNmezoMGrvBSasRujCMduNC/d+rd
OC65bzlHgtPLLgBBqtdoyeeWF45t20D7z9WdoiMCD6RbJruzWJOpMYx4kGlecgF7K1fZ/6xeMr7X
4PkrCJ7FWAbIOYo8+NLGBaEPYGe6a9nHluldDKNIAiT2d1se2Ya3iTqNq2yXCsLgyQBS8g8lT+Pe
yM2t2phkjvsccJ4updbMAAPpSuQaHTX/NCIkrl1INOKk9UJGPzTiw9V0cUIo6FZvms8qA+ZJdfaL
QuhMfGB83wg3po8oYNGzp8lIsRGOTKQN0GMFMAcCwtU15VN61LC2JnisKtDBZao4km/h4xZVUaYB
trAvGEL/MFhSXljXbHglImKS2tvbwxCwcdARjOyjDIoUc8aiEeDH0bXbXZq0xEqUC1MmSM3bfjKj
kA9rzfubn87hl61bkXeY7aGdsBGMTBhMVEqHvVvSWs4OPLkMG5WerLHLTtGrtUlAy7R7pox4ytYW
yIyWqlQFFQ0efoCOBmkQcp2n7iIYdg8+sHUQxsaPxWDpuyn1hS2N5im4U48tCG5p4pO3Vowk9gp1
V5U9PjXg1vVFKB7PWcDpiwzG54eqnp/V5yJNiM0G8fcr27ymZVvWr7Eva65ZNaYsoYHPp35KLHFU
9d7SzO53d5Qbpz3HvuKsW7fEBVTXGLUFDVC10RNrUZy4jaWnOvVG9ovthD28huph3a2PBdZXo8Bb
gYboAJ2ALfMOLIyytgOrbbMxoAIVGt2PYkMo5ZAEiOO/FPlFKIlhWFGFIS6xoX9R7IncaNBisZ4h
gqy7s12J8Sd9Aujayu2U/c8V3X2NNA1QK/JAIu0176SFLlqc74dQX/gESjw+e1GK0hdj9XIQAJ3c
1pO7qQkqsbjpr6a7WT68qhvvbY1+a9TuKeN+HnUZeGu+GDdZmTW9XxElK/FduVEi9/qfbA9CKQxO
rxcRDjZsisSXJJ7XbMja20moRdBTLxSQMv69x8mI++16eXaFhpXWgWHJrVatdWrRJRJ1JOnNZEY3
oNrujew2v1JLhnuOa9f/AWBlll0zT9DH66/Y79Ky4slKGbK54hhXxMt0aHoKnLv3mnTIxnomBFSJ
NSCGbcN7nVP8/IKfF0+K/yEnhXPNWM8iwzU9ErZwILnFq5gwuVuhV83tOBiIb1BuVP9WceF2FDwH
6V5Ed598q68spkwEw3qU3JF720QB8K/GuLKlLpja6ZRPHZMzxqVZqE78IvfQyrTmjTI8UXw6Vqvv
/fDJKEVqJwA9RwHq335gTk2EAEox5DSv1Bmmi0sQxMCK3pdh+FotI6Jbfdz/dV7shyFH8mMDGeRd
ZFoiA8KRNCNX84JFX1o3Qz2HDSknpx16B0XJSY7lZceKySFO82Yjck1ghKbpXpt6COWNZ0/7Nbjl
XX6TCVSdoiLSq4PWVCPaR7hPCLCUNU5mkunU2naBSc2vpp/rr3l0RtNAYMqKASdf2U2jL9OYBquo
Cnh/snuGgpQZFzbvAa6uHGM1Oc1yc1fhrjxnlOKYAUIXS8UOXzY7BxodaTPwTT608v4yiD7WaMPr
evsFdci0F1dqM0hRWl+ZJe0gTLqQwJ+48GPxu1duLUu+SgiU5dDfFK7+2ikDaFRApQvy4GK4A9Cu
2p0x/rgES4J1eYvoLt/krBXKDx7CWVVDws9rUN3/TUBHBPLulJISrvct/uQR55h2wiXxYcO5aaWv
NeptUCAlgZANSTj8eixk7iSniKEjH9HbyLAD8Ixq8mdKIN0wEgsCCOKRCvKJBlzQ17fyUXIAPzYt
KDxTKTt8lTrZ/+Tmw0nzjssLlyjSs9qB8KcyctbE36iTx5QAQIq4if/cT8AgtO4qCukVfoUx+cq/
hxpdaV1xzoh2N/VFuHOLqhPFje3j3pPdbJH3l0R9q3es1/7VpU3Jatkjd/bpEtBBt/cNuxcpLQco
BoGc3s7eite+GS4w6GaP1BjuSAbjuJmLqrhrm/TMoZ8/9R0St7sZvKxLGBrZvk/CYPN9tVJ8Auds
9Ti4kERi5CRRCbsH9uU1wst1cZMNcTw8GY6a7T/4MipJ8E35MtiImbEnKd/TMVPGUSJAJMhK7J7D
euj9uefiKeoI/rnxZoFLVX4lKfXpUNlLI0TbDgl7TKKWwI6THQ1LnDLKZHS3CvZRCLyMwPKH5qYr
rExETXa2SulRO5vaF7aMs/qOLsSSjJjAuZhq3Shbawj7ko2fr4ve6Y1uHZzwaFCCHh5dj+kS1BGX
JP9s4tnU11RSIw/wlNuNbd0LbukhVmz2ehZxbP/q0LphUKqPQU+nvYGwMEVzLpOpzfA2kzqHWsFw
rLxZv4t74KxV6cioYgtkn1wS5kwaFpEWwa1eJV3tscSTgyWpFKM/rB4aYO8M5Kkc4K9NhQyrptPk
gcu3WdvNj7VV8tZ/oKALt8Wjo2UE4lRrq1XYTOaCoGKDZr27baFg2T3vdrvmpnL5A4lrt/iIJfPe
9dQ8rzVYRqG8IMqWfofh8UR3pEyXtYqfU1NQYJqseyvyxf3Tj+bymlUkc38PuGJnCW0aTg72YqZZ
nCMAPPYlai6hXtIpOBRRTWeO7A+yEXLAw4uE8CCUKpCK0CFScZ9cluUGkeSfrikF0KIJ6JMgsRxL
dD2gAO3AdNOCKIPwG/PXEwPq4BuWWbMD01suqh15lzuWaK3KtqzwpbM0Ke/WYVvDcqT/2iZ9wQf6
mMsSuc1ETb75QCDcVHiSAfs7NMp1ef8TWHcCSvuNzTXPb19UPpLGHA2lAQtYY4iQ+17IrK+E/TNy
bHlbhfAMcRot4EKGnACOnvnDkVVGDYqOOsmj4FATlJbnPsaeFW6qMvy/8Rcxj8Wa8iE4P/IQflX5
ktnF9unwKPR74w9l2IP2IPIhgFGzvEyadNnOEiVUm1pS5gMOH39iR49lbWZSvnLRxLaQZJ6bTXEq
EH79GaAS5vYvyaeQWZKSdjjab2HMhY0ZKFWeG4WIuX1kzn6nwfvp/gcZety9LZTXmMnW09qiejfn
qLTsXW35tc4q/PL+VEsAqDihwZPLLfM6xx1cxeVV+MCN3J504yW56mniuFcFQmciBWymqNTRvdR1
pcbeVuT8U8xcxmf/X+qRSFnI7hoOAP8osZ0L7eaNR9zw+8syuAtCQ5DFX8A24PR7ErKHKQGE+xCj
BrY2ezShF4uvIMoqNmp9QzMCeRWsp/lWuL93+gVr3IchWMRsNtNv8Yzhrpe67sh//h8bbiY4bbWj
6OCWq4uZXaAerr5/CLNBMeqKaIIhTMjY0iTw2k2X2WpExygPH63F7KzoZnUFO2Lf42zWMZtUeiIt
Pgn9GjOCg2ESJzU8VLl886595N1j0iEsyry0q0ksL3Eq3SS9vbMkqYNeUEgKelny2CplRnOZnfj0
rdePzIaIB8bgfUERTy+6t6wSRgbCbWxYDyV+7cjcI4B1kX0bx6DkzIo9RGF86ybQtx01hjheVMFh
IXgBqoXxhYCIGGDJ9Bnqp7a6y8qxi4WYEmHOQ2SKKjFXIjGIyK6RAGcJV+CIcLCCQmXXs5ynCRuJ
VEyn0sIH0uiix3Vcnfo8O7I2eK1K5xxyuMCOijDQS3QQebNqQmUgJ28+twc7/JtA6K3gZiurbi8r
LPzdfbulcCOEpszbVTOVORDNNJ/4Pc3g9BNDrwEGhydPyMn+m8i/ex0KJwqi216OHHPExicg8u9n
SoivWAi5DrlGW1N2lUYxao17ZPKCUEF48FKYCxsWWo0g00G+kbuc3TDewMS5ZxMfDCWgzMXV7iat
u436SC9M0od4h49rQVpNq6GgnW4gzt2Nq4BirWiyg8xzsDJb24IKEm8kiXr4LSjEHQMJmr6fr6qZ
Zp9l99WNB+Be5VAq83jzYgDSn6PlwIQFP44MMMagWdjlgMQa+1nMQDF8uWWgg83xG5t+mAkbYVQz
gt4tIh1I5PA2chNeKCA5yjxx3A33Vdi5FwyhjdboyDfL0U+ozSBDpIZqTJXuvx1nPwAOWvWOpJ5n
MbRUnBbXP43Ri6L0+Xz3NVTqzcNCmU1Y9Q/6Nh9t88pnCuGhx6cbTcWDQFbr3umr4k9gkYHkMJ62
Fz4jFf5+QiYnE6yeC8l/uAW6F6UHBvp8GcGznjyqMmaygAKyp5M+SD7LZX16Mns7odGexdsxKBp2
8Hbe+Gl3x3Y9IuGAAXB/hmQ8mpl/hq74pcfvBUT4Rxt99zmXagppz64AhVj1/t0Q+ta2vctIYTzd
i/60CR0biEonMWEu58Jq3NhOK+7NkJ5PXkgVQI0UdSl6FrovhJU6S5lCuQS+/lSNNwLWduTrHl+5
5AIfJD/PCH68Gx5+XmEWwxAYI1XmHX1c8SwwpmK9bIQlFfB/uROoIfx/oqAeAGcqhEZp9qlTzpae
C0Xr9vBvxuG7RPJh10fsjx3CL/Ebeh88GP3pKaKwzw49/erRvkxAfkqAlHuFy6N+U3HFSp6qPOhy
eVWwE8PPm2AeIBxXJQ8AD6XcpMwBaVmf7fFv6ms2b3ptjKNwR6Am/NkPTyi1HHviXREzlVtIxk02
kEAVJKUISWTRXmwHVjqrhvYwDR9iF3SDMO1JNFLXx8V1TkhYPtHlQiMpPyCT6uBY6tnK1JKkLHzo
V5cHyCoTIdIcqj/yMq/w/XnEVQM7tARdkNvnZ7H7YN6+u6pkifg8MOjCyH9s6SGpedh0KUZuqT13
2msSOB0AA2QxZ4JTMqbNFFaYNb3Z9zwn1y6CYTuIU2hx+Cix7Vp6hPaLXuJi++DN3yvXt04Ugigo
VUI7ZtJC8ZkYX+dCy4ugwVtDXTUOUP/nqheZknRxJiTs1wzuB9xtN1SP/bf6PmEAHJtgQQa9zKIM
HFVKLyT7xS+/0QwaAHTUum87WI3Y8J8mbynI3zGmfTRA1KsBAAzqCH8ilVtnYBY9Rc17mSyNlLm8
1cOmhjxcNxMESNmJPj1HrMAPGBH7L3xKWNm+wzgdtjvj92KnTdoIjolzkoKTJ/4pA9PtYGTXaDMV
FaWgcg4un7Qrh2aE6dxN1piUgmksGhbO7151cNL7PAVNPvWPFEqD/oqQsZ20Ki7fUpqYmMk7ddh5
aIsVzeZE/H4HP8pnN24//uIzbaoSugo9iwr8NT9a7NboA2rWm7aay1zaqaTBUnrDUo0wfYyGn3yp
WwyWqKIbCOgAzWCgGXNJK56s5fb0GDxaKjDWo8nxhoI03/2oB/oWd7WHio18apKGbOO79t5X8IrK
X5xkR6qTuhSgh3V2I2UoWR6FUvBPI3ekPQ7kFgYh2PIfF1X2Q/dvXFO9UgcnYOlxNJUkJeyle6Rq
WFW+kJX0aEWnGagCar0V65R8f5WERh8ZXSwVVQGpP8Jtr7brWte1DPkXLBtuGqMWIgO+KWK9wUC0
xWxXncbN2uOOyeZPkXdMoszMunPoUy4gHZIPwTK8frkP7favJou75qr4MkzlwMT4Y1Fiicip7Z3l
XKfxg/DXztnwPY+c5Rt0O7V+ghwKQxwNszbxMVxBprzFHHV4cKQkbOP+iLojZN18RBhL6CIz3JAC
5rXZySijqGPK3s5vBR3MAFGkhPXx2AK9f/f6xm6PhgydnF5VpQuGhLPU1N84cXslcyRCqQZPJEj8
izRmB5ORQ1KwX+YItnOLTFRcwmXhivDIWO02ZJD+JhCyqzMXB6i1AtmwAl0UHRW5qZgqDxTaxOSE
c2mmk6/b2D5BmfnxfVbhfDznf52dwFj1sQdCAQMRaJey8exNb6lrS+0uwraYoKT9gZc+qz/2PMZ6
bssMKUasWdvDA7ylah10NOoGN5n6h016jcsz6+t9QHryhJBI7pNwNDJLrRPQUUeBHUuEKa6u3WZH
vzll5m147tNSOc7I6MWwQS9/eCBRwChlHIuAJb1eMSC9TMJcbt4E8fycN+VTK/q5PrYK4JqQz/4X
zOCouHhKHAB25irwhEkpwB26Fj3oXOlEI2b7TM3qoqiNJBvw9bn+UJ+tMbr1fP8Cungliw1VpcJT
ngUcXEapcjoY6H8wCCergN5VYnpLRkaVn9/yOx1e/GfF3Dqnrwa9iO4oL2S1TfGDaY3N1Yc9tJ4M
tEDjNhOeY8p0b65XEt+0zfcAzDJ1OOng4tbDE+RJcX2J3V+Uu7y55rKKK+qvifnNOZjGJ6RIq/8l
cd5grEiYx3B5yf3h+Bd+dc/6U/jxciQPRg5kqAnPeG1ZIPnVK9CKw0GOhS/UddJyEMl/N9fNqeB3
kywVPKC66xjuyMWOhp0Vxk6rASDCb4YnUgG5CW5XhFKINUxxJydkXY3uflxL4g/rb4dmOGpn5mTE
Lbu5b6kBbDudnCoiTb/czgQ0AnHx+fDPFZSV0c/o16ybwMBeQSDP4VbFbfSupcXmJQ1eWCyxK0lU
Ua6Pd4zr6XG707Ms4kfMbTijp2qmAf1VrrEzEI1kvHW4cH0kSjdMRHnnyq96DskyQJ+7k5OGQ4Me
sQmttE/c0/mUMuQ/9Q17R9uxCHtqRvn9scm4zXgMo/2uRYM9Iz6MvO+BPGFdC1MTRMMSuPxR+sjF
kirQTgGuvXkeLs8hWbMLHsuvw/hMZR3D+2pv1a5xE2neK3K51eB5aAjyQV9ACW8HQamiC99lhPNS
OHJWPcQRyN3Ot0lST3iWfCYxqWU/TYhE+bjw4YkplizfPoLM6ubf+uFmmNzcVLV3x+Etpv3D2Xch
S22G3+0vwvQQvjrI8CMd2Lq6qaqSuwPrnHedKWA+rQ+659Ey0+eKnPAnco7C4OUfGaW31gqfj3k9
V16wskvYr7U6HVSpo0B9/yFg7e+ln4Gqbop8z2M2tZQ1IQVyeGjB3b3lnLVE2mvJdNHalg8mcqyW
FPeicgstTdSj1H5V64tG2R19qn2PxIiguT4w3eOTHDhVwq9sLmBncvZhZNMcU1htgIfZNieVjoBS
296UFbBqkJ9uZupbKB1zHYyowBBh7jPyQxf1KYOe2NpCtzQ+xdUQWGxl/GmYne/NfnGT4kNnnHMu
6XqSyAwa5qQF6/h96gF/2P8al8VENMZnWIhBqJT499msTYmJWZ4Y1LACkCoQtEQkAAwFjYcPETih
j8Z7fsYS014j+IfdYDl56Ld6ogz0Vf14tR3IoqHb3sEz5yACPaufjgx94MfAZ/6/86b+GKJ6R2zW
yQLSoIHULDUCKz2ZQBAalmMIlSoMx478IxY3XQKTJZboc1f4QRiQpLLwn9xRQXdRaE77fIoPZcYX
SCuIBIHe7DshAOmFavdtO9bEui+qNIKb4D/XQ+1oa9eiiuUmamxhkA2NE8ikzuW0a8g8L1NBRVdC
34tfSVXz9F0zhClhI8JEAI5bwLsbTmpoyKOF9wFTDqmvYT+9Qy7U2/TBDpKWn8DNLas5V1w3cKrc
5c8Q/ND93QSlJlOGfPgiLy8eXV2DlIUUvZ+A16AUBzpBSyHHyjBgwFq07DSjX9sYLnmOPYdsUCve
E+HCW0spXzs+/RrQj2XCHcCZSJoZyi9fcicwLd147t4SS7cfVbDx+BxWtmmp+WhUXy2IyZr1VBOx
VLW/pUv5VFr0wenoAhp9RMgs/sOM+fLuVvuHy0TT/y4MmMYW7XUjJnf1a5RH7ocX4Gw8R52i3mtB
BqQLOIPh5TqHueK4YVuhdPUwbybIdUz4D0YMRW3DOirYzZWaez7asnwKW9YpA/DORLflFfW8nTYW
4lO4fGx92xo8kofiZUCF6eEjlqepXfQGuCjWoeUsRYqaEtsD7p7cgnitTzVbW67/FnJhNoZLtUaA
KPmAFDUrVGb2mJx7/rb5jiwxuCxOMCZaIU0mc25rc/bk6Rx+FqggMhxIQpBhzfhmdO46HeT7H/gI
FGPFoAvXzFSdus3GygnXdoVmN/vyQXc1eANfE1zlb/24Z4GFacbggLxDLFAkyTDc1W7+/aHyPH5i
CV+z8WOINp1Agdoevo1NDVvUEBHrq8tCW2gM/Av7NuuTO1V96N0gLC90svrgG2XOfmn0DBThZSyg
9N/V+Yu2LyuFaR8U1IF7kUtiCXTmPkIvhXjnvfXHCZnZJ0b5L9pVUwYdhH7OiWzScrlGYbIDDuGc
gyBo4V34Y8Fx81j3oI+zyTfOuSgtHgZFYad4t8Kh4gTJ0YOgVMsiidL+oCDQf+POUdqiHkECCIFM
ZNFynpn9r5eUVgvTsLE5rUvUQhkcVh8/pWxEe+hV2ocqsUZczH99uXKNhePTH54a0wvDLQp+ArcC
k2gGoFKIIpaXLu8cDKfVSXG7oIDFbvgM1/HGMyOgAePgIQHOio09wBtRP/Bfpi8f7RDVwMPvFzKn
MwDoq/NQ33PuE4tTEShygam/XHY2BljJxtMyXmPi2zxCTsjdywpi2OWKfibv0WP1UcVNYnNcSL+E
XdO0HpQGmzCQ0yey3Kj58jX6zcAh50AHelVUS25ZFPnD1TFHNw+exdWjCNPvsV9tLIPRbisKE4aF
U9xYkhLEOvHau21y60K9abqrUMytQRJ/RN1DnhvmVabK255LgxK04+8Yct8b9E0xJgjoNHYhEb5o
4BppaSZqaPlUNyYSgWX440Vr4Vrr3aMBSGx1zaWgqBtdtYsStjcmgNmYwoX0l9+N5b6sfazj0Xyp
3Q5LuonabEv1L5g98uKWHM2jE/ZN8oNGxwe9iccDLjWMNZHe1qZnOI++1U44+7pxSMtex3sZibQR
GTI803/WEgKZ084nbDUNij9tB/NcGRRxt/F6aTnpbMH5tNiYUz4zEi5DFJ7dH5KeGaOfSRBOqZ5+
n0cZGTzkjtMrePTjV2DOMlQRfueae7p5zMpWtBZf+oIfx+tjuKQQ54LeZAer0qbivY0dirKJxQOW
M0HENApSstnr5sqtmBMVh+j6WbqFciLJGvjs1cgfV8dydmuEcURKxtZaSyE5TQa1+9L+3juuzzKe
rB5HScFEuaoEYrSnj9WX2nA6a/by9zbq1TTG8bTfsvW5lAaE165Ax9sjC+XxL7ar2GqO1nBk1els
Myvia6TIQ7kkqxcSuINUPOCKMdzK89An0gXxqgCJjOxBSqIcD9cFl1VI7gYGZ59u8JmF1u33J5kd
sfWZ49sN8I3GgwMABXQYw+4L/eXeQrmhgrp9VKgDy5FfuRN3eeKo7rd7BlR0OidX4jV3rxse3OjO
CtzGacgnrG4LXdpoxL0rbKje5hvaw9kB9GVjhfZU6T30w9nWkS3J2tx3QOIvEG2LeowbLAmvJczw
Hi7ag+o1XnjiNjE2HYC3crCLN9aansotUs139DutCv60pV5IBTyjBGT19YgreexrLglJkibxzgud
sn3uNbe822fn6Lpfk1XRCO7JcnnkT81P0CWyG8lb2MmaL2RAEj2WRlveaKyN+beHex+zjdFLlov+
EUHsgr/Whuwg+BX5Zl9sMbFqDV3dGmxzoNCCPqBeq69bGw+cCYV0sieE4zTDUKFF4c+KFg6MzqAa
2L2EKAcSxk+c2d6PDb5V8vSjttvdAvrmvX/xSKTYde5RROOGHO3ysX9FZcLTwtITLWH2f/17Cdot
OZ5ShXYJCLoSUtV6RhDXHmV49SQxPJjSu735g46W+fwXuWZ555IVW9LWM4727SEg/PUpUKoSSoMF
Aoy0Kg9r2wm6YIMKiSPe4Pz0soE5UUTBsEMlivSWnHaOGXSLpKtXkiH4eWXsl+F8q2W7HwMu5/42
96cypgJyp+3rJ6KPAJkrAXtChw0r6628rpf3zTtKUtROIYz0XnbSEP8v2sxLkBw016mXokkkBgex
yZ7Fe8NBG2ry5qfp5rsbne5eUttNcEjHWzby0ZvBDo2UabqireS2qApRZXO0v+lWqDxGKyaGAod0
1VDLv/HsUfAwlbCcrK7AphCv2sl9TKuEJR576y/P0KoyBlZIYLKal+LU2P0iQWK6D6Kyz6TTMr8e
JFDMHtuXk2pvNPoh3Vpjm3h5CjSSF3EqPebS2CMV6CQUv+lxNZq6YoSH0TdnHJj9dlUbPur3WzDE
7SOtwEAwCQn1td54i9+WF5ZH9isHVkiRVfd8UNgZ0XVZQN8NRcbvEBUTwCo6ivQzBCkU+1KOsUvI
foUwxEaoAJz6cM33h5IUGNhc2lKFaMsEBEj8PVIhZBDLkM0fPHRLjVd4dUPiGj/8bGQxVtnmLD8/
7q7SlaI1FFKCnq7tu/ox6EKs15yIpH72mGKZdN6yy9PZW7rPdydS67kyrUguRpGWYyEym2WKbBgA
cqWYRdbm9qzudDYxUiloeiOxKBaVUpb8ouQ+elO34kXi/tRJiueOwIok86fDSwoWz8FaCq1x3aV8
GTnl5pCq6PEzKgBnWKgmLwwkP2ePJBA3jbfxCsso64+zYJYrHhRMjlaF9MgfXsGY2550hADL8bBK
wEsyyDbP/mDlUMayPO/nLW3QBY/d8iOLs78H1WvUICu0f9IBTwQ4Zgo0mMKGSg6uZejKEJMPJHhf
8joHadqPmjqjtTcMqu97MgQeprnvGVKtsoEhxn+nGrWW8/Gns65jPOeTPFB4NxKUEHSqa85G94Z1
WfkWjNEsmH1tmUa2Py4GeVEaCUK9qhzELuBLAXSvX+Im2SkQeoxaH0GahWlwP4Plq4Y/e0Y6UWPW
7a2fLyxJTSx6y3ivwgflvuyix9P6dImD13EPQHLtOoi2KYqnRo9wSvZ8WQ4c9N/FGlwSk5vvFMPd
/mvrjnS0RX1VsqLtiAAkT7KNVq1f2qGV6LOf+ncQ1KfmaFnWf8zAfxdBYrub9ptfNz6TqjCcJIZM
ctCxYYDgHDASzbtCA2N6X/3lfe+WQ78wsxXzFwfJsN768eSposlY9Jn9fAP+y+D3pTRRMr7G8sxn
ljvnkPjvH2qwzp03AjgXr+KmFa83phuVrP713OCUE6r2fy3ZAzvFE1RJwjjrMKqZxoWV6tGo3r6g
ubrS78yBP9NNjlMKYbazeBNUYq7UCCrXWrxrPZ/t2PLpA+GanfYxhcA5IaFnucvc7Hu51C5DPKYl
yjSA8+ziOyB0VDMOu9p3bYtLaz2ye+vuiY8vNJWFY482+AieLJGkC+j57x9R+J4nyBhTmnnSIWBI
dGkBCQCohQcUJUko5MXwTorWP9fjmhnQuHYm8k1pzhFlq2YQ65HgDJIHTSaKYcRfLhob0MbnSRQd
Q7Z+8BnbOMkeqGMW+40ZQPNh0W+rKUYREY/G0i17tAOyWevwClUGmNhR+OPTXaRvSx15t1vgz/as
c+UvITimYLWsNboRzuZkDgKB35PlxgBsLC5DpLQbXIMNHvwBtY7qoQcepAjDTQQyXeuVdxHjxkc1
PeB8JnN66VYOCpKwPNIi/1LrgiHnudzg2t0odL6VgdacVXQOLcKdtK5E2poWQM6H4ZaF1718KERQ
jM6Hbxn8/Kmif3Q7TckMmBRCO6YSerkrIKVJsqycnFQojJO99WnBu/ZGI1utOvefNUBgcP+6ZJix
gJ122KiRQlx5mBoxPGQrRfFnUXMgxlKwVR7I5IYrYJPO5PF8ZujVvlYTWnEuFMoD73hroixu2JzO
06FaabTZ1nA7b7Vadbh3MHFC0ktZ8utmD/JLnHG24yHjy28CYpUK2Tht3YWQGVMg2TSqrjpywCAE
z5JnrCxX1ORH8Rm+2grGAtbdwuvvj4RSpN7YBoPQsuLgWfoiyEj4xStF/GQP4jEXZv03fnck01C9
izA/obc8mE1PyT27zYD+niY4waYAnsMgV6NPVpWdzYbw6BtFwZUgVm47PrpObDSmMm/kwnkkeB+t
GbU4Uu4tl361ljKgZZ0Jl2q7ZjeY6EIsAh5HfrdmpGBLn1rElxjAFE3mys4fN/6ikxnCGKTUhzXw
fvodARDXoONSBJgDFOU8SaysllPr8ciL6WjqbNPmESd7EgnvxKpImkCk0VIYECUeOGvEujZ6Wn/P
IGgaCzljuHrKz7NSauHoSpRmCU0DXLL209p/qHd7idwY5++pA8JB9dFG6XlJoEBpyWgqVPUxPmzp
hCs2VzxBOyNIX1u8iuyJGWWR495uPTbqy6/PWhahX2Jc/1mU9nRO6pW3Ne9FKolJYbto0LlII317
gr2SIEEl+M7RxLsHU3ei6pMjXIlisyv4Nfs63sibqgf11BUYvyGqczmxbBXPM81zk3bCm28iTvvv
GmkXZbn2TjiEvCQZZBxtowARZlzKRU0t7oxkWh+R1Bi+VyblAtv37t/svC2Xfo5CMdzIh6m47Mf5
PI529t3EPdyrDBmGmmwhxgDn/gqtPzdXgBaHIxlJHYX3rnHZSZByXHAy3WzoAqK/9NRuotvQ5xuN
IWJZ/jfW6BzOOFH55kH2WyycbzwTQhGMe5ETLuDCx+8cfFJl4II0OrB5ZEMLI7AV5Agg321WxHJ6
Wl4hPiVGygImp3vEJfasgNv9RUK/a0SXzunaG7aFJ97lPAdcneMxWKsjtm987Zzt/6B4dPygt1BO
fgEbH0DXaxlMzQAA7TeSvZyMhJ1UcZWc3Sx1JcBiMtLgjFxvW1AQKay5icFpBlPB/SLfHvx5Zbo/
VBpq3JKMPlAg68FfuekrD/LjCGUs2AvhhZ7vakqOcJHxs5hSnRhMxqFb2lErZ54LO2COBfLLDbms
xpoxqhHcPAkqqypyz4XoyC5Q0dZoA4arO7oBESPFqYuM0ntA+KnpGf/EhCkrUOQ6nEskAYfwju8Y
YkUHPjE/AtV6SMQOBvx0qfK4lOSpCcZHtWKmH7tU4rowgs98YJNFbdDHfkWjUrqEfIDaUS25l9pH
QZxKtDbGdcjoJa7nR9FucqWDTlKNv+Aygm8kA3POL9qstA5209SH33xAdPZJWdrBpPsyj2j3p8bG
s8cQqJt7U15t4Ah29jRRNTfSJ4p5FpRlLGFN4a1HulUy68pIqTwDG5h8TghaS3juhf4XwwUF5o8p
Ra2+WRjJo/bQF/tvKm2XlNBgiso+sYW/zcZ3tDw2N18UiS2Murjy836Fy2BVx4c7de1XvxMDW1xo
51GGH3l6yu7c+BQ/BJA7URHuvAS19YuWyNbUySAO0lhgHCSRYH+Oaz4uNdCnOCmfRekyArilB3fZ
45/XP5th7gfkq8zZjUFivxyjzbCUHEHuECf9bFoWxTArIGJwxNg209Yr/E0QT6VJUuXYKZCs1cBi
dgMa9oecWahhQ+kBGyBtl1Z2WWx0x4N5BK5owlid9IILZRuyRA9E92munlWCI/tuSoySTzfMXr2L
1jCy1lsXQNSZbb5+NvUCpYovHoT+LHg+xZJrAdSDHn1Uu8R1Uh1z2Glj1uHpY7HMvz7SiBjcOKdN
SbxzGrGzrppcnxm11e7zXhKfLECYkVCo3WYHptgikfHgKEEGetqOHCEMSs3xGRu7YTOJETnAxJl6
6QkOE4PhEQZi1nDjmM0pLca66TXDAvcgO/GtJ1aiFBssvRfJU8w2zYefYG+tFWpFsU06Yq9lYsG+
2lH5ZY2Tmu/Rv5hGPCYW3hYhVj+3UixHWrkWoOGsZoKrIQ3i/krG9tvVt91WcsSzc4O1LikQFO3X
SXGTIZObYbc/RAb9Wuma2ajF6kq3AmrzxA6Q5cglHH7G00EAt/dF7LHl47dWjONgtmXkDD1PcHbi
N3rnL4TODBp6WEMVY0oQoDBy9XkKUg5ApJv0HMmt7VuHqnHBQtOhaaDTQ4c+j4C4B3YgM+PkFBES
kOPhGrS7r249GWU3kfnzWcnH+ORUmhqpehvZXprqrFCT2cPcEexo0LbMSMmtfTQlp7JtK2Mr++AE
UCjoH2iFqgcNfItjtBveVRF0JvxCDIoxwDCiJca0Hj1v+QmLf3Jwwku5sytl2s5WsRFz0Tsp9Qfe
xQCtZyW6PczZFpKjB4T3zmOMFO0InsAQZU96bR/U/NGA1oTNdwB+vvmXXtHh3MbceshVKya40JjT
fhASm3GXrJxRc/lA9zMOFO6N0+hkcZZIf+sfEzVA+xQI1NciGgI2ZxlSK7x0IAalpe4M1ZmRNMKF
hi1ckSfPAPkZicNc26+yUZPMmjgQcy4nkTBmS0oHguqlV2VFob45CDprtS6kKaGGW7NG9TdVVIVZ
Oo4qOjlY/biW9Vx58A1jyMsN9OggqnxWlAKh1Ssg+msOD91IZoje99LBc2F+6nWCSvZqe6HF8jGj
0Fg1oHQOGkRowlEflUC5gsuVWrTil1WeHprqYhTM05SOnwlf2caWw1Z5VSWwmetzFjIPxaM32MKq
+4Ke81s31iWb4kiXDBFCzGC592GVbAZFHtB/+zh4ft93+aD/Xj29Y+5QU2PgrmHVfHq3akRwrYlg
ZJbP5d1IDPmvtzhEs4uiVehNUL0TDms4S0b81MzgDazKR4M1vcjRG2+PEciKSk1UH7Y+b9b/R2Tv
JtMfGB2QnVtDip45dhxU3O4hZavAGLlUor9BGE/zRNli6I3OzR3OjmI0sNlnRwsJAE6V9j7FtDW9
uv646jReKZXTNIIVjeaI0LjvcesM0cfToVaz8YSYCWBNf/nCsoIB6fpoHHOzNK+Z/OtTegh5WFNq
C1po7D3naFHeqZZeg2oNn0Kh28xGTvzNRM9Cv8p8jG707/BI6xihjz+TYM6AXCus/C/m02cUG+DS
6K3sIwQ3Wh+1lrOdcqsS+jEl5FORcfGSCeXxYWx5Sf5VTk1EPgDdIv4YBizgWSc64gS9wYMDsWpL
38nUwO4I9sFUuQMh2NjaiFtiY+TdQPzMXhdWFYRQpZjpCWgP3F1uN5hp7CWr1MRkP6W7WmPPZt9a
WkxYWrXjagJnlIwmy93Kn+zSHA1DtQlvVwZ9x1LuobUYRVHCfsQhNDxRCnpRs/nfxDBGfZ6vg90V
2+JbyXTE2BTx5sOFYIVVG9HUbHIo9xZGtgeKg3G5LGjX/H5f8CIbJCQxaGaIKQ8vyPbvr9GCwBuv
4xe90lBMChvHjjlXBrFCsXArDPk8qR355AbPVycxn/KNioAl6DC6SRMdEBfz79zSgXwLhj66SvMT
/1SoYzVMQxL5E3P2k2EeWXfYSytCFU1E7fNI7K4aPjNqmjiDlBEjOAmzYkBTTBrLPnD4xUEOYosn
vNyke3n2WlsArPQmswn1ef4UEMQGPo2/mMXZz02ymV/yhmliH44JBKSQfbNbmYpfdmuGXSkJxUcL
sKoRGsiKgbN7E2BEt3OPun8pnQQv2vkgz1pNDkZjiOGxn7MY22H1yRUUBnUDWZrB8vzGw7vF20ja
T+rMcQuBH3cLgE6LxypIoMnxrBIJKtqxZtaOvAhXWPCf9RMF21w8t71ZP/N6p/mSJdMIyPLPCkzw
A0X7f9EwCTe+s6n9mGt++op+MGFviX9N16lONC581Mm3dmC6Ry+r2zK0rBeQWrML6MqTfgMgmCVO
1BFpdtSkGkDzLcxuP1tBtFHviPwxhexYrqr1rKX2i2hYRe3oTV8FUPOcqKMbh9pdoIwiJjygqxyB
n8BOdh655hmu8WftyTUoNCrwIrFcyhf6apjY52IiwYuAkjGShWDqypPVQZqxcWujcV+woYIsN9xy
FQiiIYirtW7fBoQvCO8mTnI5rt7pdF1A55jc0ZDBv/viXeQ713Xqz1IaIYlXsesqd3Lr91VGxwLY
ZzEp5weM77tPDuGUQ/8j2YP6r4BnTz4hIAK0w0EodzcTWb28G8dvQAVa4Q7A+A3VBt4G/dh+utCN
duAT6MnF2Vase29JW2YZDVWFzLZr0WpVG/HnwJY40MQccSh41ysM2DbOXoGE0UVCGQJEHxPdtBOy
+aI17sVYgxbGHxAxxyasMQI9+UzffIZAqZpgPJOp3Eq+1hkjCgtQO8Lm8y+idhvme7MXtcMTxXPn
MVnAzeCvI3oTeHeco0+8cAaomfIBGgOb9VbrdVLMOB31ckEW+FNsKNnwr7Nkm6kfOi5ZMppbZ7G7
EqaD1sWkABaz5AEL4rzSYrfeh0Bw0K5YNAMcstHEKpGtKXm1GFgF+RMPmhoEkjwvAaw+8QFhJw9U
WsEpyWfdOYcfL3RuwA0VKhZk8TjMSJ+bOs0bZu9+8YGuk/fcNukFNJ+3hqe53JWkSFDcflHBRvFm
0a0Hm5umuDnavo8WvRGj7C8aVlK5TV3pNcmVdJYLhCZ2lm3HXmQqmwavrTZfQCVBlzEBFLhfeLuC
qpI8QkRklNWqzsxdKUyWp+Us+MocBBg6yLO3DPS8LuC3i3MUDd26LXWXoCXfCq26EoO6vK90ZoBG
FsCt8DW/WuvNXOe889ZmEeRfahrtmrgQu0c/KF3kHD3a9pqZzWfl6UYFrRUDRROJiLnkRACZJd6q
bktp87Ic4m52Gkx1q5JtHZFpxrmgosDYeSaOWl7+iUIRdws9wMS5btR4/qrdhZLKKX1RVnX3BBCm
4/2iehPXg4u45SY7rupLjQEj8Z6fbIv8tOr28wc7m9/bFX5mKwfODpGviMTlHZpjHoBtCnl0sjaE
SHVbvSu3R+3iaZMtd+CCgTriOEDH0IgbrxRyAVW8wBxMlfKeXqvyKmSk4qd/poVSPyqzbiSsNmTM
ZbbosSihR7LisBbPEWy/y8fUc9g55vWxMgJlAwRTgVwRu8vNL1ICmDyYXkWOhgILLsQJq9+EagQo
JSOECfj712Ebjnp2lrOr1KWvmnrf9M6vSzkLeJUKoLgmpkjDMg8DGJ3QeH2nL4+7xS1t+Ipd6+zZ
iucUWNHAjs7P9KClsFA+KSXJpFbF1rnM7lzG2IRfPbaqXZl7PT2ZD1L5itTlT92eC1yQOVvRuJad
ew7aYasywhq63unpxMeavW4qw37dxopLjCHzn6rJ2AfVGO/ysKjD/9OpMV8izDg6NdNURiMdhNTo
sFOTorKLhsHe+0QAlA223fXqNzR0LeJ6BPjPRocGEwemcmbm5DoFWiGOTJhrVhVKkFvk7WWHoS0e
0qTuAsc7YOHNIq4YWwJh5UsZH32TuN7K3GsnyMAHxHIhSHOfXqwOJQX83XQDx+f10s4a0QYPrja0
dcETBDNdN+gt1hTUDbu44AR0KiHTgiXpaJqZztk8jZvmsudfb7IpGTACPaxQcrkykJh0OjdSe2th
sD6XsjG4t7C/rdc7pqpqF3bEuAcH6vSDB8hXIeXik0lKAOknu9tXq8ndTRabIi4cDNim5c7HbgMf
BVRniPtUOFrpUJNuCCpdFG898D2sWgn7fXP0XgLAKAoQIvKkg9GKp2h+mA6pXLrYtgafUBepb1jY
jrcSjh7BX8vGukpGmsQmxn8QvTpKDrbMjE4VL0NvETWIq4ZKevw72ibu8A4G/Myx7siNSxdrwq2C
PDfkne0Cq5doeH6BtNWcVbgJs83QU9T+gw+HPzenno8hA0YTvH87vjcGTLQuaX1Nzfyl72FneGzJ
RJNUOr5+V/KKOUJyOeLjzoGUXmQ5OURBXPEvZ/h1TpT0FnZFHv/SSyf8ieyC8t7X+i/drWOeEU6i
+5v48IC/PDRECPK/leE5uxyqledOfpAeV3IPvWeNEE+huuJEvZ5b8y1Dlg8WwIiWvjinV4LP8Tja
vx1n8DygQB8fVpO9kFx4ActB78OfUwVLriYhTLwXMN9JenEDV/oMxrD8MxUMdsjYJNQ381vWMacD
1+iIfngfZLp3HeJ8hqJE8ZC/JL5388O0mKQhX1sL+L+o3lkVd1ic45N46H01Vfr2ydBkjXo/5x4V
wkDmtBiHz3ifyjKSSXEYbjWbzHVFFIjkLrf9JR0GHivYcFQt/SwJyc1RZa7xBCYKy1doNCukV76u
dv6BzR+76YYB3M0sHM1BIHs+WAp+lXIq1SHvbwLfEkaeUCrMFRvF5tHiCzACVyej+969E1oGyDnx
BMHq1wMdxc/JtHf2mRQa0lSELHdba+632roK03pvcIA1mlt+gtBsv9JbPhtcB88BpZIcOubR0VPY
zyTyfgFnmB3TYF6eS2uOf/583JU+92y9B3nDLKhJzLKz3rKoCYygS73d7q352zKgGt9UxiVCA4Xz
QgMKZk92GukXoV/3yzr4gl2ZuhywpB6FVBdaoo31oqYTK4oXhlqm/AJgk9JMwcsPJ+tjjdrY0LC5
ozUUhLN5gIe0FqGBeZ5JltacH+ODvthwiUGkorDxH3V2fdRFpjqlBZTsJ2duP4ID8eG/3QntaFVA
Tg77RSsqoTxYRyfqjY4bEsWyqlCVkBe5G4xXtJR5z900Q/zvX8d2BT0LDh+6vRMLiR+WcgXKGd4i
gTMEcBJSU5LD9ohydLoYCknYqEMju1DFrqtuJ8s8VWG78bR6huVkmBoID81rVRHGnbnMm16Gvscx
sVtV+r6vbLv4WEAxG6bwkSPag3t2/dbuWc1a5ZgBb2QqyqvbC0/+64J1KKfkq4G7eqsS1XqbVv7G
I2j1lv69al//rE7NBmnnIkbZKT2dRLh29GDFB4cBVkQnTS8HGDIjCvpYsJHR20QlJnxpy8/A+VKG
qc3jrMBLadvn1p2ftoqUe2ekbjoTdxErVZ2uM/izL+RC9x9CQJmJOGQaHCiDilJr24VhEgSD1qnR
yQGP+nZTHJOBZL0o4ecji8MXuTJy9GRNf2hTJOOMEzmfH9hDAZA7HdiZ+kfFPvF8dUeTS15zNRgK
RWFDFAimH0Y6+YXr6OPyHSjVGl+Qt/EQUo3RzSEdTowpK/gZnaZIwir/cqzZ7i/lGY1mEEoI4Sar
o24HvIRopBDUdh/qOHzVyK/yKg/CuRF99LusiDsFZh4K1Lg6XaGOU5pTEJfXfct+qrAR1uQ/nzuP
fFvRvFISJvCrkNLcJTYAIhCdYZccocdF5fNVArLumgfTRFLpa3do3dg4IGWJ5RsNVKo5O9STi7c1
c92oA7OnG+K7n8IQCT6+xq8BPs92PSqh1YvpFRaZ46qzmTqofrwTkxz3QAIb9/omXx/3kBE6u17Y
MxnYVWfCpAgrJ1tEbIO/7VK+IM/pdxN6lUvd6EsQ/sUe40cSskcn4hpPUD4g/x+CJBAjEjg4zOSD
S0JARY3U3zLItcK5mDjv9fCP0hbI3UzfjaT7PDukSYKP9LrskeFqVZr7bxo3x7sUzhnIWCWzUhBA
aREFT3c1yKALRkD1kkpUNRcIPKfnfNOV+l+fSgzMKNlRE1o7/s8ab3uF71cXIQtLQVsbdlhrGXVx
77OqbadKlTdQT8dfkJqGjzMQsxkI/j2qvxVWA8D2qE9O9tvKK+glrxotFCdi9ACVLLQuLbnhdBK2
FEpWD+uhhb4NDVndWjcPfs+9lvQnyWNJO0ocTZqNMv9QTxgqsB+7FreY0VB/ysSQusoQVY9fEzON
6vt+Vx0UxRZJEbuyhxufiHnjVd6NgumJVlMb+N23fCV2DvdGgLVW99yhLDE0eM9OKAp5TXj/V4b6
QbV9XIqymxVnC3U7cHOTb2FhTBwrQ8hp7zuGoyHUuum5IZUiWJQzs8KVZpFH0QaRJ6OgvuriFZTt
ReaLpnPrY0ymiDgj/lAiu/RUIDZO4ne4jX8IAKHea5m55H5NwVgiMkBeuAwN8NAvnbrcfC/IHGEV
uZCGC4F3LnCTg2MY/KZydv8fVoSqBI1bZrIT1lFN7UE8Sr2dHdNdLKq8S2g0htt0NmpiGmAI5Y0h
N2YHXSJgb6TYzDIQSfAFKh9rHVJvyCsPr1Qt/vrbaaLU51Yy1XIDeGswetIVR0zJTiTn07aSXwt0
j3O4utUrQltpoM5tMrcjN2pqMmWeU1mO5sfxCCuF/kZdowjkXnt6tHP9M1sZctROGI2StuQHXGYj
tLzmjt5ycKy+RUazwC/aZ5KzbkR4iH2jFL0jO/ONohReiIc5UcuE2ElPxFiM+GBm3bJRV21l+5W9
lhLkagHdo4yH+y1n6VC43C3n/QnxHYichKkve8wiNqH7jnqhFiYjCM1VsHiFmYIoWzKHYCG1RdIS
kBKtWD3fqwMuRp04/t6dUp8Utgn0dhOeNByDN0NnBxjmEcvQQxAkl3gKuEj+FTNnuM7lyEllf9YZ
GuTijGo8sDzNGbYzxJZuhNe+0ZMGu7xophWlMA2CFWFI3+3025dvMfmSv9XTvNVoFFZkF4KfMBPk
urDIInxyoJiaGwHCzLmswsNQVkeymLGAaCLjyhthFnGzogvlhLnxTjW+rl/uwEViZfs+Q1eag7EU
Yotp+FqN5mmAy7xKu9TJyDVNf+kWZhEPj0fPtoB5w6xLYEjIDs9HXsbkYZI2ph8utsqLiZI1iqqN
C/iVA9WJBqwg8cr2A1jrGWy34xvxo2A4WZFED229BSumRJPE45ZS7flTypM6hEVxrOLyNUS/SBKM
aj29WYvVAwvctRJEUKO4rqLeU6k17vMUqOt2ylboNkrq3hXdzh+YK3cR2Uo1GDOy/iqxK4lADZ8O
WcvxhpVui6Pdq4yA5RbnRQTnJ0pNvJ6U3XjM/0ZUqXciKoaT02LJKryOlN14bTgUkGaWMcGZksSR
wGT9QbaBqc/+14t4yJLAMk2Cvk5m74blcWKSurRqrbAFMcy+eXi+t1Jf8QqjRhHctrOADj3LQ4y9
cK2EcXapNpAD56vVjDetMW0OefOI6UboCR4338Rp/9EKNAWMH+gTRB//BS7kBVEmY90VOAuUTiCW
ZnfOTqi5D2N4KBFTLcQe4uoaxqEsqi4GvUUpj5M0fOGMUqbYIqXLiDoi4nJ+peLtG27iQHQWqJaO
roukmAZq1N8NmAkZdsm0yHgGsNjMHqNvavMHD+bgDz2pH5d0MsYaJqu/lFi7639+zaAp8eF4iNoy
8Mu7rIdPMnwcFLOfTj9AlFx7VIoUUU2Hx1WaebBC2ca8ohjAHb5ay49HLuu4cnsfRHqcLijSne+/
VoPcccBhlZpf+gH4YkxTOYK4H95jVOn/KAxNUNAhegNT65W7j0NMj9KseJ6J6zPvSLXBguUrs69+
y6hXXO+jrpq//Xmvj5TNhq9JbWnBuEOy5yW9kPxPPrLux6geCpyOtQ06pjKdw86zt1W1UltEXvQJ
28GTaTSbw2+qixAyRTichW7JyZFVV+lXVwQSKVk6lI9vtfK5xIq+EMqnhmhI33FbuiJwv7Zs7uf0
X+cjszXicWvp4GxHP5T57fh7s1LPEteAkz2bJtCVlnDA2uQv/26qnZW+3T3iDVgTeoGnVwo0jpkR
Vf3NeZm/EgCdaj9E4b8z7x98bhIzdTw4e73HCJnyd7qvtep4mZoEzXFmmjoC4LDDuxTx/t7pX0QM
Slwkr4kJFt2IGU0BynAzOcvJ8Ry4Tm1MQBrElCq3s9c9ViUgNuBrQS8AbmkGSmgHHzBe2+R2z/OB
3wfBr1QrIKaC+yLP6DgOAb5lc3oQjbgZa1gpu31A6Ln5/BUcuQApZX/lFzKAFiqlT6vywKqP6Tzd
bX0CzVb/qBxvp3c/IQ46BbXfnabOzAFEEzeEjS0EXtrA6nPqETGO0QQ1p0wjtQqtVRt27Y/ofjuN
qjSWFG3actmtN3fkEbkEqwkeI9P04N16zyJjT8ROkMHOw9JLlc805FUezn4dUB3dYCtxF+vlsk19
Cwo2boeHBCidNS3IXRUI3ydqp3mOlO+zBad02dq1qJkDlW0AynkS5CQzS0EAq3t/P2cgkGUGKPt8
EEk4s7FqbtemK+9cB3xRq2dxkZ8vEsfNgwHr8y1bzO3OY/MtDPLPEaSeh4QOqWt2Rb53Fkb2qZlW
lKm6OAYMlIVXr6uzZVr9P4GoNymB2MQozu9FdAOFmzjbSraowmtNXYf0kYpLHWB4+inHsl2fJjhy
FBfq7PzTjNZ7+UQLNfMWT/vyygeND8GBIjEJmYAixOnYJ1qAYRCDDJ0MLEkaov/rn2gJ+z6vsF4o
DTQjBLWns6+Dm71/Q/DEdPvP8bdO0WHUFTmWjnPOR6V8Tz08XsStUOkMOBIfYswy+9jcP/1DHw6a
MqXl6DUjXHGxVgyKQ4y1L1HN1Usik15FPvHvWoHJVGoeFjorjpY7eRSNo1Ys3LjvrUXqbkydrvX9
PW5MIfE+y7VDqgBbWIm+wyY3alZttncybvmgk2YFwoLwytRnaldvZWGcgZRXf3I3vg0L/35Q6720
Kf62HJPZ/PpbjrWZv/v5GN0UsslY+8QzYO4Co6bMcX9bn0yMEIZqyBpanctfRIqMQ3Y/Na5XdRo7
A7BuXPh0lH73dR0UzjV0kpVHCcOwmoi5TynxKcsLOGlPWGw34XL82orhpPcfiKcQ2LSpdotahM8k
nf7BA62f6QvU6q2f+Gl6LW2AGuZ/1T5ms/zHFGgu9l0VNk2BqtVClPCoaWZAawBLNSQrc3Os/HXD
czR+tzJ6dJKx3Inlmauae8YMgvn+ymSaqwlTe/Jwqd8YeqTBtGwXYsJO5esZMBFHj3ebM9cXN+so
Oc3FteLEwDQiVsview0TvEiOSnKgqdIrZuCNQlhl1PCYc076XbaJPAsPVuL034llDtov71FbgjQ/
DGj8NA6/fL0lh/JQp9w6PbcHLO8CjjqLNyZcl6GmzUgc+vgswtUB9sMwnech/SBcq39WSmmOygHB
xFk4lTjKEj8ugnO6WUgytT/2nXchGeSKwpDB4qksgZVG8uSKjUD+2lRCFkpV80YN536HaLUgRniK
Dmhz3dC3yeEfrKny9GRna7k4H9pEVJ/EJeQpCehik2rfzgMTyERUxHX2n9q6t6c+4ilV67/IsPkm
Le1/PWGu4nZ7pkzVFqIcu/X1IBXawesvuDwvuNMAxYIIqNorWT8usEve6QIBME7R0HDdc3flIjF6
mGihaj6Q4PW430h6lks5KKMZN8iK2m8lCe9K17SQwa6wB7ZqmLXfMpvu+SQYMN7DzifYAar/xMQx
kSQDWxVJp8gmFU9+8UnirB8Ji77jfkVQEpn+uDNA/P3OzP4NNaz8xWOKjaCYwoLdmLpneAmJ3jRx
QsRfT8h9Wd3Zn+dUWdIL2qcKGtYTP3A0Q/wXpJRS7Bj9udOX/MBYYYy1r2ipzkZB5ntpQjAIKMPM
zC5bmyjnL+VJSITPxxcxd8dSPw94O+a4Ws4d3uy/Hg9FUioV4JUQIJl4LhswQnEu6BAbD7RI4LAM
NkRm8gemSsh1M2RBxuscDADU/KaV3PTVEkXfK1kM1ExaCWiTEJRXiDXNcKcghOeg1uTRD1gxkggo
fq5RhByoSFnD+2/ErcgDPnZztvfEvfENpBpB8jV6QEW/Vh0KD63fGwBmLWI5lKn8k1xw5RINM7c3
OwF4z48XLla/IwfL+aqSRXwyptwOKmrWGbUhyCc/sDHk+hima5Enf5OIFenGKy77YYmhghygRwQ5
vZO1XuWk4x6eIxy94BXyojEuQy4oJjXKk3El59IZio1b4jlpzXH48Dt0yA0vYkM8FXWHsjRHZ8Jw
XxZvm+f2SWUn6+pEqGaWBDT1R66z8gE9JyJDh7O1GlsBck0dth6KB+E4ste8OUfBI6mW8m2ZGsBj
kXvRG0sQWd4Didiv9kxtogGlfywKcJuYmUQ5qtI6ZdWsJ1ZjI2ugjictBunH6P39EEF5ta5i+v8X
CPCXLx+z/ZWdyJFoj/ZfjSGV3CuTLxecWifykxeTosyIp78XUAeTtj6XnR8VRu4wDpvVkQmun2tE
/aXYMVU3RsSPFYFgzYSd2FlnzudROeMrU66CeSwsD5tCLPVI6KggUNvwbqvFVqwXEhdm9d1WG703
jPQwoVGO5C5FwCXRBCnhyyMlOSWASPmLj5/bfkAB3NVJXP8Vjh69ATAd0zbWpbogIKtyqggdJ52o
/+zDHAj9hKyjsKEVWM5BpXY78qvBHft1MgUgeGohKz3TyeWc+0Qj15zJS/vQ/WwaHw804Drp0+Br
CwAGNQZjPBsn2crFdqAaZpk7VIBLk8cUhLvYGTTlbijBbXRxWhdhjRDhw6/NslSA60HJq/SaGdfY
rOSBYGNDe/H0RSkLo0u+9SfyHLcVRHzhGliPMVmGr2Up47cW95a0bRjQeIYL0kfxOAPDs4xzV2mb
FQW5b7tef/dFGfj5mtAaSKDBqmW6gbWsvFw4oqds8mGQD/Lg3bM7kqJsI+ExaIaT8ytQeG3gXASD
JPjYsBuHH2d7MiQAo/bz/xx2B6zldHkLj9xcMchdUKxFZCcORN0g4FC5gDjDCvf+aQ2YQP7fLfqk
PUlEOT3H72HScKDQPVy0odgnY9MilNRrPGq3YY/PNJSENdgg4nVSDDOZ4v2d+BmZFmV2v5USiRg2
GUy7U1koX4br00XzpMUnA2da+iui/Pva+z0BCIIBNRYOSqQt8DMymyVefVB2DnehA84ywm4vRkN9
h3CdHSABEkOA5t/TqVRfLqHBrNZh5umqxGLuM+XJT+IUnzdx0Qz5Kjn2rrYqehIxxSCu8+Se9UFN
4sEKSJavCAEPvrHThOZN7HTgFp2166qsXBmO+YNteRkDC3/WyB+OlGiSEUOKv3iS17nK/7ylZhaP
vTZw4mwS2Dena+VVSIi5satHBTNpdp7wN02CSlpPwBLTI6BZaEOCi3TYn8O/jvf0eWLjnqNdZyoJ
mYSNncaRt76pwunvc7Guel71wXok86MPT04R1lnmdHkXaSYPULJAdvVIqb7qlRYYQQvo/upKNl4E
rWZdJmXd4rrpuCYGsnVSPfZMPDGoXQk/68J65aQwcNaWiVS2AXX5Da6MkDti49RgtrMmkSit6vi8
wcs5XraHw9N3cmShl8YJwS/+52qTm8xKQJOK9qDCRkaIXiywSTuEtoT0onMYDKz96dAFIymD9ttJ
NBJj4V3xogc2PkUAkqhRxFVhkXGUht879a9+YPD6krEzu///Rnihx6Rz++5a0bF4W3mq2P3WgwlS
YN8PSaPhqzCpGG6eJWjT/LL1d9HHGdjL3d2PSE+4jmMQqTHVg/q3XKmiTJo06phm4nW3RCql8bUC
G8ojYGIENYVQstiZiN+OUlodgpjtp3InE9KrKBpu0YKOeSWBVyeY6SoHGbRfMRgHmOZQK+Zp1qRj
kQI+0SPWLK7Cq9/y87qW+aRQcFzl3A7FC30ZSJpPu7f1IvyInkpiWh68uw1IIxAIE0kESSXSjHwJ
p4zKbojz3yyvqVX7oYnRDlRfQUjhbudqlQgjhQXrJxjHDpX7BS9w31o2T7w6gxhGQ4EnCQK9Z1ew
b1fazlG8UuGv58dsqxq7YYu37PN0Ypzx3F0IJ8E6kzDIKDbqQ79Wg6D7vgBlORS13rSjLMU2qEe4
RDgXjuUgCRFeLy5UXBYC8+AsgWR6H2DMBWUQ0C+rOI+1GZ7THJnPDwqYqzKJU2nU+1RBIjkQ+tyh
3UHf2YOwJM/5OMMqpYipBcNX90ozHjlg0rh0LI67DX670NfRn/0GyQegUopZyZ4hJ9PFdueO1RHQ
3UqXSoBj5eLx5w6kRQoEgU9X1Wcr8uamRa812/CzCSkihAMJktH+txKQrsbChm41mJQ5PRzP4brc
TWejWKkyNP85rZuDyXP0AE3ACg6tyz4x5KZcoDYDI0vGmVafnvQCS2a+tffJGIomGmi/Ud/lTw1R
kpfaJDW4mzSiuHcd0r73cmaZO8X4Mw7dsh7eQLHslJJnpL7To2/oueiymEY+l4RwO7nWDDkhnGvZ
4pQRo3dxfK+GD06aNs4MtBunNkBZDW4U09zuP8C086zk+5J8Va/02E3efL202a7ukhQBw3XwMpkQ
9TYPFkMteZJUmXQQDdyeEAW8Qqp6xvWQxQ/Tf+CikU5ZWnaTOm/u/X6T6pLprWInZhlZ83RVshfq
o3rpzyGYfXcWdnapwUdrsmtF1QKxa7qsW9TynhYUg9zKINZ3d/IdjS9QjlkWzEykt9RY27blAbCs
7dgY0Jd8bj4EbcJfSN+9Vp+/wOQo7s2NEhSHYX3As+D55kU9d2stTWgC2htZJMrImxOh4RD5GIoF
CQdyU2wb+fmRgcE3W726WF0w19tiuPUc4sN58RthapbyQ1F6NGSEjcfTcHP7Q92rZYlYYDMxgSE0
CiMxPKeHKBMBYojU9bPHL7KAXNiK5zLAFTRKGomz2EcKxY+Q8J1DapwCinEtjyWRAqv4NUYON1ZB
QckxfaqUtUd80TYA2knmGC/x+AFAfuGUaEY9PAlgdFzKugx/xfnA0iGQz7RTnJ3BKk+HfMp4elfI
Pby31GJAWNxH7+6lmyYbl+btcuRjuYadYaTXNu4409EF3TkmSjRYFjkqNX56dMCZfH7G8rwZgzgn
i1JqFUxgSJ4YEn8MeXwJIMDRy8NAJAz7a5DkLriC3eBv6Hyzg78S5Id73bnTJ1Bd/DRqq9fA8ntL
5CH5Qxx7vOHboF3GHqr6eD6L6ujCHyu8t8CHAcUO2SaWQcD4wGcuOlXL1i3orIL/Az8RwLtIg+LV
ZPfCnWRHfoz7432YmaLUNRGwG17yUNXgqxA7GVBGAjE3rmVtIPkccR7m3koKox4U4BnCTmho/Hth
nol87FI/tGGUQsea4JDp6ZuIT223bVlNs0FxQS9qUXB1IxT/c2z20+/YGUpA4MJ8xjrJaM+NzEjy
nIDNECVUlwR+cuybrOTgaseb3rmC/XCUVCH+vr4eV3GrwTXWr8PfeCY9jmQSaFXcf/RSmU0atFfa
DbbRRJf+7fFB2pFklU5i/VyI/AB0YlfGo4nf/IV0EQniH5dii5CA47OP5x+RUAIL3ukZWliHmFKf
VeHUQm+gJ9U+CWJVzEv1zPpuSVdWbzl5UzBl7w+U+V08elRbAelR922Y+myO86kMZ67+z5NlBbnH
29FQtEvoPYi66xiUha7U/Jg0vGg2bJEwCzXnuEh5Z+/58C0/3vu6/OSyYoVpBNqiRWqvJpub+WMv
46INBz3vdH4ZYb8yYwZyVwNMG6UY9dp6o/v9ByfOjefIvubiIFckEryLY4cjoKFNM9hR29iyl/Le
6udBpZsKHPyBU+H4WkeHWi9Le74XSi6oyZO0MJCYeP0hJunfrzqsTdA1zVj4GftNWsgviEdlmpXj
gus0GAX5iKcmsSviFvwCEmbB9MN4IKJapgW7qImgYAoC7/B2g29PCufMglkd3Z9qCbn5gLAl7qIs
mAXXaZl1thZDCy8pV2THSO8B4r3acUnjDQQ8wXTFBEyBlFqbFd3YzWJft+ggVGAvuVsmJ3NVyAYl
8Tpnkw7mLyhKz3JO9/J7v+h0PnPGjWNqIA04TlrVQzA24gvLzoTWrfKaLVEyTdIMd/opaKqqP0kv
AuoTpsbopZNoQdrWcb9rUZR1iQ9wd2CftcACYLSSrI10knHKtQT9XnkA2k2ssudzGVDOrxayMVr1
ccXpcPZhSREjSXjar+xlWA0opHsCHwZLgT8GzfyB/1/4aN3XiWdZ1WeRHBlDnfh7kP7NRUG0rlO9
1FIsxCi2eOScLSNpLgbpDAR2iVIbcsJoAAI7aLwfFSOlCVyyNOxFZn1AnZXs6ehms/kiVohw0Ath
JIjs5FqiWcWw9mdzMfGxNS7FRf38lXDmWuQuof69GjIlFTRyFgQdQUbIS7LZzsCxqS6dd2Fwj8SK
AY+DGKvQnzW4S4rIR+xSusPirodT+cQ60wGZStWOs69/GUTnyVfZX9q5Xo/EFvrf/o2D5+G3FhKP
9BPYhkwYJWm6atoiNnJmZzLhKDpH8dhfmIT86kFjABHBoIvlsZ5sYJL3DAqYsItoxS7rmTaKGD06
WWqJIPMmB3dLb+YmPvNIyoL2EkU4mEgr/HuYNeQyXKwlKVPHAr8dPOs/qpqu53PE31UNlFJyK9S2
7UAAF8JmqtP22Br95qiYAORy0gXKBX3q4jLG6hyGV/F9l2YdkQgWESnjOaT1ziGTtDoxeHR2N/r1
XQ7W+h9S4OuviCzNeqxfbpgY0kmtqHVSaccoZ81pY+FI9bjruHmtOnoQTmqKZJeAU4/Hap08Lzrp
IyM7mCmYPYbTozK2yGrSlB0JQCfPwjp9dc404iFD3T0yD5DvJg7mIhplwjkgVGzCa1C3fLsvrr3k
zXocaKNy5+PLvu2vd+2WO8sPfC4sPw0EoAgfAAtvv/vT7EbQB3LJ3NWiuqK9pgMXzgOyU39AA+Ul
0+0j1UZHCqYuOg0sMPn17NP1U47ILcz8eBa26GjsAJrxb923eVRkLim494BKN8E6rRVaJklerLkT
kN9AO3W/32Skrcq5HjozgP5438FnhR5gdLt7f303BgkNyW9/EZgyuph8B6mgoDpEUuvuYRNDOscg
0wxrB1QJz83aCgNpz1yQZJTpnain6O/ce8E0CeelR0/Azat141WCCA2FwR9GBrtVbYgwL+PvqZ6+
gff7BjeTugVTVUK21spk/gGOib6OgDiQLP8I25T7k+qGWBozi5+G8lg36g8qV0Qv1sMu54R67jKK
+UN7VmO7yridffiGEwdSbtaAwjEa/IzyBK+elNdVrqwWe0hkQUS4WZf0baY4Yj6Ce5eIWGKupcKa
ckckbl58Qc2s+1yXf6z7AGpIoAc2tM/hL6DJYCcCLoFLvl5F3oTwOkiO5oCcaOMdU937VcLk4Ljh
9RkDFfjTkWgOlTvxrp+YM10rWhxXSHL9iu+WufVUt6b+kgi785JpGXkk7+xe3Q6U4NUrXMdfW0tg
KZVMi0y7YnD4EIxax3Jz2sN2BHBQkjdpdTc0ReE/ddUxjbpSnHlpSNzbvI3Aafh/DheXSA+c1+eV
zCZ0Hjt0lZJByDFADcQi5vEaGfNPbMwlTxvo1ebI4Lkbop0+6x2RvykCCdBrA9AzS/5GnLxv+bLD
4KsLic9PXsyOcjsklzrMZkGL9Q8BrZK8kBwJro1COZ/z5ntlUOFyVmreq1ZECYD/pK393znmBdoK
CJcc4GaxDOsPLHLVbbXV+qFljYAr7aoGplJpg5SjhSYS1XGvLAXfXcFZdDOpqTo2xtC5lU05+n1S
Fhm/BrVX7lKTDjaQDOfVAesPFFuqyc2m2mFFUUZw8YFLMnXq6SXIBSPyF4BYQ2vrNCrfXOMPmhAr
QL1TpPWN2bQeT/wgll7Xg170WJmkTc20BXrU6/G8lKkyQx6qTtLYu21S7cpJMaO0nrGp7tGiTER8
LCW0pwzGHv3FBfUwDP6Gu0nLgk4Vl1+2ShHPnPQK0XCKKijrDDbQv9EbMtet/3ye3ucWxpvT1rxf
Bua/cBIQN4WNzef9yL8fxWf/J0O+DclyQ+jBxss774f5KrEUy6g+QwtlZ2NilbGPMCiHRHaTdDt8
H9Frt9s8JCbGYWcmCLfjYmB23Tf6XUCjCc02AM1rUUD0XdIPjZNukfuCc5GPAzbtoeZfq2s0jIS5
krVlhzw3ASCnvCDUec485Hhyb8h+kXdsSGLqiqFf8aA2x1cGtxStng9iUMsjgUiZbcUO9cNvVgZe
E21E2r7TdX+jqGoYo6GaTYYmYCRFJeMdB2UwBM+i73SLt404kCHaxPAk2SZ3rAbw/OQUd7ZtEBnZ
bHxI7RqCk9cJohm0/pF9hx1mKCAIShNIfW23z24jYHhyajamzQhDH/9NGBjJSKhYCGkwsndrbao6
0h4kDLLpCuOsQ4vcgFxMXzDzHTOt2ym7hgB4zw23EBI207/VyvaZXf6P5HWyiv97kcKkGPabt/Gx
8hUxpxc1y6C0r6+TrP3UR7Oi6RcFuViekvoKgk3T+5fTYS6KBCAy+YZ7wQlLIfG1g5n+DCTMcCOH
X5n9RGEpAyk08bZw86w104WeInQ1cmx+9A4+HFKNqpDTPdebvj1GdP7F+mUNGwMMcGxljTcFla31
e05E2IEwnDuyw4vhDT0UguE4PbJ8q2tiZQnYUTvzsInI5EjaEjh4sCQqjXKmjbMlyeq2IoqPfJuM
p68yG3P3pmZIC96OuUFhJHfR/3rQdGRhMfTWKdP9zWYelgMhLkkyKmQg+7ZnYrmgvseStq0KkwAS
GxNQsIienLmqzWd9kKHs6OHWzmscezUxpcZfyTvk5vIfYuXoZ0bgW7YExCv+Br6Q8uJk3VM2vT63
MLB1j9oi/o18QBPQGkJspUvq9hqUq++HudeJ4a2pojioBCjEihFg2yHJd4nrfRASuU+iZGwTGG/M
UYh85GEtvqOp9SFJfBTBga4Fvoj2IAnRjVg+wgmfCm0F2YmiZn/3xqRFt38e5gm24pFsd+eS+qZi
b29ufJPjAw+lid2FMCBh/1Z82e5bojv/Hqid9oMG8DKR2sxfreiQD2Mefek4gTNTv1oe6obCbwNn
K65ZKAoimnNaMVmx4GCdzx1/KtIQJgBsnSQKg+jhrB7REOu7Wjz43Stu703js4NGRYvIVM2Sv7fT
dad8o9eysJLGs9Ej4tjR1caZ5pmtnUdGm6m4DY+kpGt1Q2QdV0dwIR+SPQT+T5WWU3Mb9GorcrpR
EmmKJqLKJPaYWGs3rGA9pYrx1jbGnMuRzvOPCPqvW6aVdGlHN/zg7005ifcRVu+N+U29AHsIPCuJ
BbyGHlN9wMcVWcfc4PYErkwVPM0uDEoMtzMKXfDwqPpw4c+0wmAC5TGKVQibsB4xUPuUC6xig6w4
/4t+uUTGbgMu8P0YOdbmymqAAYnMP+GUCbZz9TuoYaVksaIqFVNeBKXfut8lhaNZNFl0LeHY4LNi
aKkbmzTzcHZDT/TTypFcduQlXCkJHYF10T053L+YW7eYvoSDTQD7AiAdE7SYQdUB7p6CfDQtGg+2
S2xR+FmWemlJDz83kdytI1nb121jsWeuRVmoWg88f3lHzANqFYrdiYfCvlTWeEWPZhxsvlTiafXU
03yjzDyjs4gWdI5nrAwE7tmJMlVWw96O8rklNAyRWW7gIOGQx6m3N29PFknspYdxmdyOgT3dylRM
0KvROhwU5KZTXGW9JyTnRyCRQFFqpyznxUh/wvzZpF8UGtY8Bs38XRAOkb63gi+4y08JtqFT7Fco
2mY9QMjZ58wtzGoCqogB5FEd4la9mrD0fL1M2UQBPyklqcxUP7rBtZcZhhPTZVFlozsZjLU0kq02
JrmCclmhkMbpJZRVKfiFRFsV1ajKAxOzegNSWXf98obQQqySP82FTqYU01JePYcAOkAh8Z9EP1Pa
/gx2ciEiPB6yg9kKoTA61FcOtYnpxMb5cqMmshnIPS0BoAU4x5Cl5SGFskW3ihWj36Fwt9hnO2ld
2UFVuWE5fih/bexRs5b27md2bsAbotSq2JSgK9PVcQ5YF6LSZQgDSYs5CS40q69V3jfC29RohXe5
bX8MmWz05mleNEiydbLAkNDJLnFrkaRtYIw8WvXhiRXYZvVsx6CS95k+RTzkEPXh+nwcbPMy9vAC
AQG1YSH50eB8AWZ/CycmczbHNcrdjLIcFvKmM8k1f10oIFvHVBHq22HfiIwAP5MO8t7CNuwA4xul
IvVhomJ40dJoiqZJvzGMKdNo3zms0oJzjjEcpdHh9N1Y4zl4pogEtKCsUbGf5WiUkZ2wkntuwVeI
Oc5EFIsPQYfpzgIMPl+NEj7FrW7NIThNn4XNNBfuPfHgkS5wRETqwJT641y8KkkyIrXIcl+N0CIA
huaGidP96eg5VQqlAEatlvL2wElsXhrcSzAjnakiQ1tpxHiAYL95XxakDGmK3wNJsW3pz0ICHdFs
Xt6AEiolfdAX54ru2fehq76z5VSN43LqiOAOMv/SbpCXTAxvEDAy4Zfjdr9Qrp83hpugQf7nKP7W
Ihv9tmTCL6Xe1unihT61Zfu51nvBbjNmNclsuzAMWg87SoUAnbB6YFtsBvoNsbyuH8b1lhHTtth+
fJdGuB3Lgrxl7U/0T8ELg51chNxsLC3fF+2N2T8ZYZ/3IM5rJ2WlSt+BL11OL3Sx5gDwNXubG4tR
aIaPtmsIydaE50C2TYGEezRq5zDFCFGwg3+FN/2DyvIWtoXCyHtDUMVcm3ptZGqGc2m4EulGgEXx
q9odHKQx10sblcsCGy2liuakVXKvHFvku8mwaqn7GOdSd/gvXIJ4Itmp+2DrNHeaXuoFqTb2X4DG
Tn5PKKWinep7oD82Bu/Q5mCH8f1QW1YBKp5rIAWe76XiVaCeR4CtayzlRYP1LDCSMfaJ9Vp8hmKY
a5WtbomxfVp6+OnQfGKQtkyT/OX/00xQluiDHH6CaMCc72qodp08Dfz2QeNlX0jv49jOWtipYuF2
kQVb+RCHxNYc0qjHSVGb/djfa49y/bWGhFx6C8IxWo8JMjKH8NaNJfM5BVU1PNQczdUAW6MuCAPY
U55esUu1sz5xpISLwL8/EKBpiqFZctQGWaeBF1fR6vEG6aZcORaEtjlEFiEur+hb4FDlM6sPN4vv
Hnhl+pgT5TOuNFsiMzBqBGYhAISiQXs8sw74gCjE7qoqWU5SRestkEON++PX7n/ptCoKETaaSSvz
s1p20XCpjlBBNJ+tneEoGMdGw7hgE56e9vmzJhaAXlo1OjIGYpslHpsh+HiS91IikvEQjVz7SqFy
CKX1p7w3/py7+65vzNIL7GU0aJmb9Sfw/1UrcsbRw7HKojF1icE/N3qcZzBfZ0wkFutBFfx5kQX3
ydKyG9T8GcGBz5xD02LR8qWmdl7IBvGokhQA2RGjFqIK9TmY0idt807H2dlJRrzWS0lLZ/0kBXhG
ntf+qN+9T52zaxrp4cshRk8QEzgQVjXr7Gx6issRHVHnC8bJxZquBacyDpCPEp31RBSOqRe9TDXn
N2KxTnERsVc29m1xrmRq24GGfKWEK/BAuVmlIY2wNEPTXm5xIbFe9DBE8W0x5qghG+kQAZ587Liz
++/9R/JzeqEAsWLo95hxsrx5A34lnWCBwHD7uQHPuLyBc9E5OH7L02CiZoJhTJfb+MmRMnlV6qJP
V38bHgUU3qMPOMNen/obihttG3mx3EpQrHOy6K8qWAtKnyuBzcX6HBStpLRwlFe3eJiVOy9WjLYe
hjk+Y3hy7KpSW9moiYqe8IaGHNiZgjXgdk0b06uzzTnZJXj0HEVC1KN4OSA7uIM2eGm0zEumSFhD
wgUbfOWRNZt8EwsbEZ/JY+BoPNuXUI1awH4cyAeuFb5o8O1TF723u9XQinZNouscywWneSHqjqE7
3inUyoejz+G47d7ENEz2POfyA3HHh+7qOh+OjcZgd0DEf8EKOi9sbsP6ZWkkV0jrOdF2RM6htTf3
pHYJcydNZ/DyLSSd40Vq2mZiQTflYDzddpcWeo+6kzCCEtoFjpom1ATwvyk9ZLgFiCzA55KSZJkT
lPzin4TPos0sPQhbv7eGc9T2XhB2lmb0XZLNp1YOdwdJmi/7twA8dBWEGGhp8n2THMo1tp51kWWS
UIiy949on32eVsU2HdmnNVNFwOv8glzAT5VPd7RXi759wqxUtb2gcMHm35RxWD4CmI0LjcNythcp
4Nwsa85HIc7B0M8/OGBvqnfPSOJXy7ZezESTWH9Q2PDKEUOEo+tXJqoJ1PFPzNSkxJgR4WcnXeg8
nC/rxM6lW3GZlsOvJgH0+U9c/uimj0/Ez7WHJ4IwT7nstQIy2BwWsZ7DObS0or9pY1+5/C13rVLE
Dz8JvSgJe50sOvQXtatxv6xeBAca0MyVxWhkd0dQvCWwufR1NATLudD9zKIXkX3pOVyDvAO4bnGB
o/y13iInuNPaC82BR3dDKtJu4ZP1LDivN309M2lft1OVNWd8pUDirZzQXKLCkWu0LY4nxQim8m9s
NVLlpr2Jx0xS2JLXtIKFN+RJA0fNRWO00qqPRnRQXNW62EEC+RbqfG9Ag4muzxJSL0WvGAsjbZZ8
6JFZxlaHJ6DtaFrE6pBi6+HnjyLtji9OhqKsZ8abRfAnjx2dERgrVr0LtRt5ZiqyXks/KGb5YV4F
hE701hAnE0hPmjVI2DPV1iq9M95wndBxTGH2osImX0kQ0G5ahYWs20MT8utuqlaIO4LwVbW0cYca
zOPBdYpePA5VS3xaiW062rRbTD1HmSXLmngHFlWfYz+117sJCCzPYowm9TIgE+4gpMlVajaB1fTr
UMEw2caLoPtgAuPNbvSGbwXCY3Y1Dl0VaWHbXN1jXtcTsd9C+Ji/rN6hobBLbrgnZBShj+lxVoC9
zf/SiuEsOZIapUkgN9dKa36sBc8Mvdf+2wlaCO6FJoMDSlnpaBGX91OUm4CSwE+lVJInPqotzDnK
m+qG6PbwZexut44Q7g1A/CTd9ioQcOiSABnhLiS6U4Os7Y7Kox0384TrRzXHtQol2SvR9ujc+AWH
phoF6VGcRanU9hw56lcfejU/WbL6rXHHb7+R+biFKyFbY/+0QxB3jejYh5hfCg18cUqk7LeZ9A8g
Iv36GJhOFaGTUdLu626Bjum7thU1MLKuZmcjrJLoMVJYAJapA4xu4BWMnKhFaJNfx0BpJPPyDHq4
C6fv4Yia8kmq2qMm/Vou/M9LzQ6pPgpqCBmDrD+3759rzOQh1isjlHv4uUgvhRdH0JpvGw0Z6kkT
1o1IoJMr/MlRiHtotooP29dlZ+qipNNMGkdiGf3gcWj3yIu7tscxr8uuiErZkhQuPJ/q6VUMg5Tl
cGqaUJn+05/Av0XhI6htGFoZd83/yFwkGkAIMlOWi4Eg133t/L2//hsua0LlT/VDfJhucO4b+EqA
YaU0/m2c66WNOtxUMLx+FF3UN5dbRWrJMyolUj8TZMppNEuOU5gCDJV3IkAZp/XlhdnVr4U0LWiu
YrssJFy218lq9sEPVMlRnFwoWB/RodYCcV+jBnFyjZ2bsXBXrx3lL+1V3vBFNslwsvQhlYLi07HG
Zm/aSWlC1KCIJfYItFm64DpY7ME7g3DKGSgKJ7WwKafwocMxh5jav9V5yTweaopB7P17rdY5U4+D
v0YTBp72mc8SrDgwVj1ssDqHn3Yg2JYGL+QnC2+J44rZ0o08BH8LYd33Iqq/mY/AMlg0P8zoDaPI
y5W6CKpYLW7uQQj+UaLAHmpbjTzO9cdg101r9hsmusPNKA7QuY2TJKPrWOWOvm0E7/U2eU3q+XD4
JwaCoi24yIBPZuryqEn2bQIKhfk0yP8dPGl3PJAojLKvqhYHZaY+xYDfT7lHgzcA4gv0eXGVquuP
FxX8xg6lWZf1Tn8bt2I4cnNNpnZTfaq/MkbKpaO3ZguNKeS59cbx1QRd/rEGelPaEjXxoTrMn2VJ
ya+lgjq5Q7N9Cyeb50GCvSZ52epVtvX85JX+6GuUkI2KQNcc5u0D9UidEsGZMRR5vxYAFwZDZsOw
poblkaRW3cKV7SM3PYYmlIiNPQAR6duQWT/LBXAsJOGL1T+umGowoJcnDslRSwy13U9Bk2a96ibm
hKXzCZ0+MZEGSaxUq10L91jfm8wFAGMoUHpmSX4WIzAKF3P9oEwwxbdFVjDL5bMHfwJYGR+Azogx
BlM+P5sBvK5Qas5TcrW4odf9dIXKe1BzCQIMJ7ajh4f7AJ/+Oth/62SuiHyjlGN71GzqXWrLWhah
C9G6Ifb1hX9NzsCruGA/vHXmYZaabaetkXiAPSUz/sc9YZx390/RsZ2uOt5d1qcc1bS5R50IIyeD
0AIoIovvMt1Wt0QT0ppcXaOWdbVW+baydb8Rghu6+plzJgGQyuqkUzPOg7Q9taGk9FkekQh4YqKZ
PE65CCIkqSDo7L090AtmQkmkYNfh2DsuIFV3GHZQWQubAresH+Fm4i7fRrlpPA0U8KLnhoKhItCS
SciVbGH24WMUivxLi6qjTM+pJOSkao4njAs7tOqkXLOFNMp2+4e6vRXskWyBPRAhyTZ8ENcaNwJw
UOdvtqdeOe3xFDtQrDrtP1dB3V+TVvJiegS2sBobtwmdSM5dVIRJm8V+udO92zQvwXqpaqz7i9+P
9koqTE44R5KFzHhzIXr1VyucGdWpmpo5nla6JmmRsw/YG4vTkKnCIomo0H8P3MA1n14/sPtwKdeS
Hyuer7UUVri/nWrWzLkL+NhEnGC2xckNXoSgSYHLIEu+F5nJpvz6WnnpJc7smlSLDDeMVbal3SUI
FlS6tLclsRWb9GpGDYl/bXCAGwjfi4zsji1vyBjPeLzV7LnOc4Ep80OxKe/5B6vbT03WyK195SNe
oEZ9hDh8M4U9nXAmlyIBGoZiupPydeUJhcrkUNeDLLMutA775zagAshDSNe423ppJa9en6AAXPqb
4yRAP4D9G/w6N06y19yDWmCJrElRtIMlbZLlsdo/wkdDjKGPC4C0tmhacylqi6sm+kHKnwHZr+Qz
xwdwWWYrH+t9s6WyC7sW7HyimlZDFhH1oiYMrx3/mssPH0sv/nGQPD67bYcaWQQF+t3HI4bazQis
sESRqkZW9iFc57rcal5MsbCJ4KWb7UpleaLDwFxvoC5x46T3F8wlx3WpcrcFILTZN+pTrD6APxdD
N2mHjDMRHRU6uZv4RgJWfmBAU9xQyIn2MLxDkh325wzRizw3Njx9r2kBbTayJyYpHvICXhK2Hi/t
Z9d1CJOSL3uDgcDOqZZstq8umBAZI1x0ew6TuZQF+Fba6EuXB7alPgDQTm21jaOJM/hLYlyuV3Ja
AQrYx2GuNNIqx8uESz86n2XCsJPeTnS9SebV41+ye7lBM5f8cW3VGchqA4XyyzQxVx8X/XbvHZ4h
tRv5KOmqWl07OnKrmI2jlouahGHjg3GgF9jLauOor5c3X1ztL8X37FbQXNUo3kNwbPLStJEIW9r0
S6KpFAZorVXKY4gUQKSTADqnDbNsWvgcA1eetWTWOzJmOWn9IoyhtTuqYjc1901+ujlqmCRSq6bk
lBlRD1jyWmeUjKf0VSPRJEWmkxEmmCnDu2yAHEQsdEY4lxtXABVmZv2K79TYz8uiH26CP8V3GgqZ
J9bSTJ2P0gjDomDtzGD0tGM1D4e6Q5nEjyWXrGx4792HveOFAri2KWP3cAGcPV/TneQVY7fC+ySg
QXWinKsHEEomovak+CfZOfBOU9I1qaghjN776AGoOqcXr0xKegwTaTW0JvsHlJyMPNjJrttjyedJ
XYjQdOdhqrN/Zy+mtR9UHpM/3jvUgkvb3gEWkQ/PUtPext21F8LHnTn+L56zMQUymlMkvm9HQvVT
S8vvX90U2x/wDa0pFZXd/r4kx+HDSvKOb/oaG5wCMUcVsV7IvzseadwbI2PXYtPLiuqUUC8KIvsF
Ladwqf0+xitczeAKQHIOKi0jr7OuEdO+u3ewdGqHyAHauk3X4Lt3hsz2IQtniX19OauaIbOYSELf
aPjEqe5VgihtL+Xj/6Qr2Ge6KzhlB60MTC47hrU9CHQMQrVX/Oj32LAVsVLAufdctiVx/gQJ72O9
Jth6f2oSHXzvqZeW195CHKPydK2ObfP3YB9wf/J4M/RJWbP1aFRHGQKzGnVpd36tPt17zUTLV4G+
NN1TUWYz7b+xGnudizHzBoTDXG+m1+KmxAYgVed9WCFn35Z+iJBIDaMRos/s7HYd6lgMBAH6nXpB
ZJZCMALPQuSZE/GRypJPzNNOPZ+BXwWrwKEhr1BXlmNxjAN46N38EXSf8dYbmWyEgxSpeSwBCUe+
OXdDsqGgiQU7M1erO0/YI5tWVRjyILeIYkC+wdutVrbToR1m0nqK7FIt/nu08E6fxLLPX7MCGIIc
PU6gJRltbRd7hYGdVcrhJxrkzFC6I0iILVV3c1nMzzHYBZ2S/nlC95qFZYIPaVgvJfMJwiGptrlY
ga5czFoBdq/KfKJ+BtLquJRiyCWTu5gTiQ64KkWHVJpe+xsEbN85ZB+eTV2xE00e9tVcnsYlJRLv
OQqS1hGfbZcOsFDaGV0OOFlbcWmc7zOZ/a4nlZOCQImTzdvOLidZI/G06LdOITSVEWbhgfisc9dr
M+ZWRzILt8X60ah5GaPSocuwYPFD1jjhwX8fJ/g07XGYRk+5Fr/BYRgNyVMgBl9bLDfXuhOq1eVM
EFMQvOECOZ9/a0CjkOVZicqlpl6QmOsyHBQA+9e98ZAVyMPAz4QKT8ozoJ5hnbgWYDDdajLMPl2G
Il6/qw1swhjdms9R4HypFDZS8l9i6wLQ9GhR/jM26F8gMUEGMHKF8f0HUCtEMEf6VXl2wPKaPIl3
qTLs4O29rL5z5sOfsYmwN9npjEDEWqS3TqWqK0qhk/v+G6lBjhPi+POBxia+sKFhaXFVpYmCW2n5
cti/gNnwjDBoxj3MzSvIXpIjjAymLYzDlBmAPPAOCVLXkr4XlCqMRuq/UWIyqkTQ5Twso1lT1W77
+nDxCaozNz+J8J5KqktNafNu1aJVQu1nR7u1VFXndBI29oDQIYNvHo4wJVy68ZVpwgTeY0Fs/Myv
huYVs8zUnlFhw32mLlHuiZ9uzYbY1SJDlBE8A21tV98exZMLkveH59TLi7/MlHUHzFzK+PWA7nGZ
QzFnwF7qyjcdxWbBRoTOZtDTHXHhRmS9f1oQPvvcqwQ2h2JURjFqjvXDdQha00cidNYM1nKnQQvr
FIAaLJg15NwZV/lXQ7GEpckWi5YpXJ6zMfLjkOTQdDZKJdImnUh1PlVeLE+xPsxHSoKX1ke4O7+t
u0Bc6UUbN8TnzGnct2Z4Try9B2Clt5scXwP+i7IXz5LP8bYC26TLXDrdxvYNZDeUZx9ensqTAugj
e28NlYUvRGylCknehTnWpIYj1oX2ItYuU+O1LpvdweXo9jzd3amgGLAPYwhV2NVdR9dNGoMVuPQF
rz3Uj9F3Yp8lgPWsOwVrX3XzGFXYmtAydjUe4tWLY/S7ug0J3NptDnD78AtXyFRsdIfROEjfc0oM
GSJkRunz+IO5Cj9R/VpuxYLisb5OhXHLDUEYts4XDkrRouSLyJylPsx9wluC0302+DV7jil/G5xq
KOfBd6AJBWQbeWnLnfH74f2ob7/OSwLUIt+XhHrT8hPAyj22HrspY0XT2ki/J+3+h58a/Qgboz7Y
jz9Wf6G00mF0YRhHZDOXnaCzi0qvLkk0U9HU79SBumaYP594rnTZC2/bTpNUVzxCgGSWCz2/ZJX9
/2Pwp2hUmH5wFN5GCf0aCXui2rhLIPHY0TGyoSRDAY0EC20b/B9wtNB7Ma5d74Gqgx2KsGSK+NuQ
dxDYVdwV39pC8sfdbWV3vGVlVPfsK9qtMwgCop1sHIAYQacX1wTy040MH5VZdRgR8RKzCOpmNgfx
dwNUpQVfUZPeAqSfkp6ZfUkXp1K3s9fp0Od/KwN2sGkJwEBhlGsylv74h8Uff6m9AJqQ+skoSBYy
dlLAk2qosX6zKXtxt2ZEuqr8D5JbCV73pe3D0aXow5PBpL0NBvUDUqxW1wTWl3rCPaOfbN80vB70
qG19GjQSAx3w0ZX66OuhyIC9Q2pYdK659p6wIm1aXIf2+OO01ZMDS2bCo2VI4MATC2tdBLMJDEGX
181pLLnlJFEJzp29nUdNadFsqmEQ6VVwzMzGAvNxS6k/3OuHS9ox8mC82UPUntq+bOXl00BWbSeB
QUoXuNKvUzZSefYBRHc8waJcLFKT2+HfDmJuP6Zn53DfIefws3vF7GW5fXKRQWNF3vLnmMMmNNwt
3JI+NuP9gFyLhNBvR0Vji2FNiAEdJbk3WKIVFd6Nir4cuWweSghcZFP56/4C8sYB+XMrVpd4zBzt
J5/WEd1AIxFeD9z7aoucZa+xjBa8wpnE4+Yo7jiNY5p9Iv5y4p3+kitEIPgMjRjAgLORry8llsiO
JvRnZedR6JRslpy3rHLWYap5EvTzZ+gu5bmvToxfWu0ewpCpgJvqMEDcR2fyFeBcy4gJ5RecnyjB
bvVAy2ucIvFcZI19CzStjk1DVKKpCey3qVv+HEJ1XqynvLOq5MdBrqpWhVp8BKvriDzveMfzSSno
+YaLVlsYkYvIgI5sfVh29HEwa70IsbFyj3KFP2ennSkaStNtbQy+0VlZFbePVLd9/u2HR0kldPfI
y0lo5+kPM8QkI3fYGk1WwrDjzXWXOPDPXXjB74fres20LlnY0OXP2ZXDkyhMEiyO1cZ95h2sCKG/
8gf03zRPL4UAptjMF0aPsUfWcwTUP0j+Q5ZAg7x64NTc3GCgfMc8eh6wMqahpeJNWuKFzpSBbG1L
OUkNwZOM/ay50ZvQ5XElLjm6xlXzO4NgQVvOdBcVAGEB1dZmoyHCC/lJvACiEjo+AMy0jrbOVksl
GHf0+KC1gi/xb9k2gOrvT6ZmMwQ2Ba2M4dEjeWPmgjIzysQ8xeESauPMBpIY6Om8UwouBqA8OLXp
RADdWUVQ8PAdaCRF0+vf+tXImz8o7hnaoYENkeCBpdgnLjs8HQVyk5wty8VlK52aIcqNHi56VnZ3
haJCy+fOMuK3epVEKrnlimDbxhcpK4IYdS24J7qHpsPtiFzEYc2IdJjX81l/NKR0NdEfNUqIhxYE
SXGxSaVa5NrxuqMSEjkaGsryQQ9YrXWCVrtgEUqoWshUdAm2AXXPJMEWyLLHnnimzLMhbi7if+jx
S6najpHtZC91Ffpj9j7jJ41cTYfUDADip7AaaI1jMakoTnOrvZav0NgN3w2tjBXpLsy2MN2CaEi+
eSR+vyjB/NOp6PGZPnZekO1h3g/QCXB7CWdHouB15dOPYnz9LVXg05aWYTMFofQkdG43Ue2sWeQu
hqDjP7YSnc418YisJTs5g0yrlzT3GC4l57hJmC/wRJXWd1mfneojRZJwhCQaz6a7etQBcsYVmhIq
KsbiZwJe7+snNghWk1XAWuY4XjOthbrqLOwWqvi0C8mveUzSawyjDHiKDgA529V6LPIB7IXyftkD
eyxfqQal+TGpt2iUogQ2K/sGi5IIyboyZXOW1FVxA2MuxwHsAYYHBE3XooQdtniMY2yX28FOuhtk
D54/Rdo+RsQquS/mnENVOnCoOUDuJCf4q82bRjl9WGgVycsitYvH/Od69j/33m/c3SLTuoEXhRcA
jShD1ttmv2UojqLHe9RaIOwwoulTlGBDswmEAKWAPwGW2DsNWpKFz/zBRidXMt4y4TCexZGxWs7M
KWkl7TBScGHddO1kC0tg50TO7LEQFhMQSaVORDThYYUUSqR7HS8ip40lj/CCLfNONCkiWTzOeTqD
IXujLEZb+uX5MoudFt7wdFEgNKcIgnWNyZU2jQfzCsKDHHJ6qIHRzCiSK0szWKRQ6tgv685vyt4H
hJmFSb7YuBBpPdU0TU2qEUW3P6RWEu0/kP1WthaoIXkJ8+d9ELoAHNy7h176fe9hOciB4h3Kr9tI
Hbxq4BdHPsk9MuY3PY8Ggm67sVcHSI/CSM+FyO7bfoL59jnU4oZHlx5wJXJZ22TOa9xXEv8ohnkB
yhOGLnW0/geOhB5odiPBcj9YJMr2cOoKSN/UyG3U3ZzfTPXowGDjYsRrjNQ+qOErKWJm4FUvuN4c
U1XA/182Z3Of8NDjOEbrfhY7aDEgNeQOuPhv7LWR0LUSaBg5Jo2rcyqwss4s5qx+aI1EfF8xLk2A
4I5xyB2YjT6C1yHx9I1p6pSOxA7k5MBqgGUH3OQQ2W9dHLRc/TfZBMG1avxrUwtiGxFMrkIE8+6o
hzthK8FxuMUXMzeL1kR4Cfp8cEUOL55E1Qi4Yox6q25cbjgu9y18lKkcMS9zunGLUByLOz7iRPrJ
/yB7F+vN1Fdj+Dl9qW+rm8PqDx/Aj/kZQVyKLxfYng8B1qb/yQvaGMp9y8vgqXupmBhUqlbQ7dfe
DhZc9+l5CxTFkA9J2CuAvOS/BrHU2atTvHNLTLjzQIoHS3BQovEIJ8VHnS1DU0f7jZVBgAAnJ3jD
QkJ9Rhji0AFK1eydj1VTfNw2llqzzIsEIse0G5DykKD4QjAqrKVkEB6afAxGZkC36UDmhRG675a0
svbqzj/bATQzLMPj6G45FVZzh2nSQQ2sCSEW/sUN3Eu3t5VitTt0Zn1ZdTpq1px6/aT9WSljZNzm
UVCrpeSzJtDPCB+ir7dttqBuAdbA7mgQ24ofRqoLkh3s8RqvUgSYP/dYNpEJEZlm08vTz4LT5V45
E1lcu+epVy2mK6XTgLnc2Zd2sedvPE3cOgDukDH1cIiiLJ5F8qA1Zt8atB5T7wWYI3uYOnP7D0FI
vEdHSszyetD9ewfq2h+eCOL2+6/NNHmzKtfX3264HXRuZGA7pP160j95dHVVc44v8Be3l1oFCuN9
QqSc+talpwF6/ZmQwKBfGFXkX4bndxGagpxWRyLQt2QHNovkbwuWtbAORF4INXUTTPj2HvbJf6Sd
YVM4oKohFsXp/S6QfP+KeNRspkD8vdCmGYID8Huzd1YkNZ/WQRwhzJACnRbpEbcQ9EYgwRGXf2db
b2Xyb+kEM4+GVCXEp5+gwlcYQcP5yzuSKZJxkSzG2dPgE4EqzQRAClUa7W3/EZXUnbzllS1hL8KW
kRrzssoPRZV9iiYpKbXtz0NidaDE/7cqB6BMb70cdU3zxDw9LdJLJVrffMgo9qJbKkeYpTheKjao
Sxs8wzpEvRB1GN7BM5gYiAHG08d6BlrXnZLS3T5PWLpKFIetG7AUxvWMmrSp9ztRcsTs3S0+z/c1
t3n8JMpsLxdkk39FRMwOGYYO7azRpzT947gNEm0nJZaOufBzvRqy5gWjiYt1gqHsjOB0BdRowRL4
pZugtpNgFaetlP2mb/vY5+YyLqe8Zpi3lm2NalWd0VPgw1kfsAr2IburjKGzzntr2S7trsUc4Avm
OuVt788IF/1KfwPqf3Ju+LWguwgWk42z2DZLBZRHHnqRG85JQrwAMy54gaIL48B5H6FJQEiE009s
53dr7cr6Ta9D0vkcyUnPr2IobuFbM3AgmT7nVoWGaVEOkrjIuOs6cwKiXFGqyWjX+0vYUdZQmUXk
58NnQyvrbP18HevvSGgRIfXavRT7p6iAduNmWgiwdojYwLhxszRHfbS5FpcTveqnhH/13Sbz2kCv
jsmNqq0ORKZo7wDtTo96J+hwS3y6pcs6e3t9I7f2O+RfN9GNOjQRlsAX4JI28II/m1UK+Gg8Pc67
o3QLHHBsDgUYCWxNvbcOLO1reUoDxpWxK6yqtKp7LEwz6CWBXn6SZZwXXR1bSRqK3kuYNIe+k28M
yY+KD9rXeZLD2giep7ffaudet95kec+16+ax+sbEkOLPHd9KXX5O65n1DXZOdrBq/mnVGmrSIPa2
9TSR7+BtIzMq7gcQ0OmPEu8aSK3yj5emhFdniFXcu6P+zzQgG0HxnsewgcY3yXFZ41nhfhLn86Hs
97lK8ar6wPqQeuSaaFkTuNpbPVDbiGEVwkZWEVVebhr39m8vCoonkU52DmeIhGR9hLCCSAY04eC8
CHDETwRL3Y3JaY/+XUzn7tpK18Bt93ZIqXBu1qSZQqesa4Sgs0ATjlQUtueq7PcmYiZt3PfULT3b
dHQHpx/fKmDyy5JAq1E/0vDw42FLyHOejwyFLuSix/o6xgTqQJFx81W69u91RVHToOceRSxTTijP
WCrHWvbhUAMz2my8V2Ds4wjidjkAAbw+szZ26XcyiaxINLBVH0gx8kwfdjn7kIhtMY6Ny0RI/8iZ
ZKOYz3RL/SFkXvWvKCJ2InQTIdyY9fr+WdwX6N1e88gIYwQPokclkq4T2IJUP6cvtLF1GuKFRHjL
jOzmyMtSotEvJJXoCLeyr3mzAGwXnnhbhVkfTkm8JiqjkAXLu0T9LeW8zSgLyrCxOEu0LYjzpodv
LWT0XHMCC2MmoUNAOPK59CwGybIak3LsuK5WW2JHivVHmQDgl36jYDIZ0GS7Mcth6+Y3HvCwK8Xl
DhZ3i6ywKJltX6B4z2h2mSnMPrckA6uYiP1bshIhiJzF9wQmw35BysSTeVlfNRj1qq4aHXzA48DE
sgtx6qRAxiB6/O8nI1ppmG/v080K5FYJo9i0Vvovdl3OZXZyc+C0UrHq3v2iiShNZxNlo7IrLeCP
vcLNkcDvyG2cwLoSmZqKfYT6OJiDMkJBgI88VgR8iV//a1LyLSh97rXoNo9DOSFwXKmKUzOw6Zch
Ad4zHCyzLoI6Zxs21jI4sOgbMTIRX74zlRehjqxi5/n8FXbCNpiXOvUyK77qcld0ta/ifp6Qk1Mj
QEAp2Fl2eKlX9Uce4mmfJFpNbn/mDA3f+3eD0vVTOnpUWzwRj+vf607/OTfvZTd6kmvCs8LpPa3H
pQAOdakrTsUPk4jMn4y9kTDXVVE6R9JqtkepU11I+0qzRDchvMtFmYDSLbvexDN/qYdeSbIZv1hw
IEm/eG+wBGPtb8vsGkxbOLOJD56pLgeHsv00A3spsWHZvx3Z+kjZAPG5kAWSsi3jTv95fltQ80nh
3LacBrvWgux9fJ5YMAVn99BikTyCvE2ChxhoeZvfoDqQeqKw8ZLkdXVegmOcQe8AUjmKQ7hNDV7J
uOX9dCd8TuVsHAVydBVfGoBJDLaPW7egAvCBzjnCNJecyTzsDzEumjB5m03p9qFvy02c2fnQnY4P
TbQxke6DuL8UOWXTvNSkC3FPXhEgXZpZbvQH13cg1xBcLXnsOz9Vqar413K7YDp7SwRy4Jvs+Owj
3V2Z0+Qq2OtRxa9rmbDehNyiewFk5zpiICW3HQ51okpl3UfpygBtQCqqX/4HaN/dMhHAYhklXVGq
62XRkclkFez+OK0f5TIUnBcQ9ktye6TRUo9hJNpJjs7hKtr6KsNOjocHe+7SJrLwVZ3rAA05bPQw
+E7NH5NIeMhZezitkBW3/j7TIzFb0Tb2LzXTDbpuDC81mGz9uzs2aXtHlro2/DwkGRfEm+dIKJfX
nDzMKHViMoGjg67r3r88UGs5W7GlZ6dM3CQ4kDRJOL0CpZ2GiC0R+U8TRrdwcRPcpj+lENJSlXVT
rqNP0ClYqDfUiZKdYNC/zpbmqTPy/yeaBkN0vli5HheBg0p3U74T27/+2SdGDBq4SfSHP8HkYESJ
Uukf7/hRrPDSljxUSFwHWzvVRYx9xF/nxewkLhepOBjlaE6OW5KuRYf4bljzggW90dJiyPvd7TtG
X9IeMiMObDXNyRKp+DM9l50ZL06Oigp84/xnKc2p6shed9++HDs0W7jWhF/0Kz4/1shnvkaPnJBe
BpqfxzsVu4PFkomBolPOxdYftcqMetWdMFKNgN9Fh0f0h1ju5ypOB0zedYEM1h6vx+r1jtOkhtPI
SQk2Kxl9OsbzdeF0Sa6vcY0VLJj8DUJCvsmWF0oN3Qj2UV/OtBCA82Z0ywgDfuc6xJhm5VeSK745
t5f8eZhmSSZQXIfe2fxgvVVnfNGHd8H1kePwAlpe2RqheVzFRFMxuHF4UAOr/a3eR13P0BpXSz2l
tL44unXCdvt+I6QhuNaq76yYvNXKQ3PfCpwFxZUYTqEM0pJ4nH2nz7mWdK046gg3S3PTT/8KGtOq
QCmmVEY8/DtFYJjc6gDz9JiVNYK/mDjVWKxvu6FMFWg73Y3vK4hmJzufROSCch2n7ZhWWTZFPY83
DFjXoqjA3qzQE3csqpA0/JaX8KLD1X8UNVDaciQBG9dERVEGA0lWOPHfT0UH2ICjSnjyxXAPN+yU
yKklLrGN1tJNV8i5Ely2IhDERUcAgl4qBZHWjqkWHDd1s1yo2XVaEBcmzgeQEh5LFU+lP3m/0TKE
a6Hev2clxpiIM0XYNYkJQIhyHOn/TqWCYL/Jk0Nli0teyqHeP207Bt+KzABQ5U+Naug4/1B4UXQW
XBTBuRhjccrosUvHdKEpwo+KrpqWZuuT1EEKsfDmtsQs9JqpdzFoWL2ppUWEmRYVd/QCZZtRf0um
Bpm1v1SmhUi+KiKy17SupPRNxJ1j87CSyclmfKEaUHbHWZPK3heOvWBec9uRMwWJmbsChOHUdEUw
PkJlyu3O+cldak9E5nhXUz+9npQKgkqSzbAyP+/+x2/hkC5X0SJB+mFMnYt2utPN0ckGxaJQuDzx
NjJGLF9tr/j9iLqyXo/C0rUJTCrGFiJCjReRhHoDLsxVAFMCPJnQJywpzJssGeq4SGBQGKuv1F7o
vVS/rlG1uxqT7CLS5VwV2pvOMc6B86eK6hW7gUtAOnFKRDOM6hjc5eJ3FUwA9JVk3xAPBIGXC7Xu
WjVkpxTy0aC8Q0HjZO1Mh022P7UGtRr9ys4SPOHXgRM/RypbFTskNcwPXLv8D9JTGgDhrEYWnUq0
QJoDu2QZzqaoRL0Y7JeF2zqY/+agLnjBQex+DCQWz3QCj49K+qxHrYQ2uYk9DDoDyxgkDKgMPo35
+g9WBdGICa4m7ATbVaGJySLewPDFoSWYd3MFjS69FBBGeRLKcMnvmwOfAKli8INT3fqwjeDQX9y8
80OBwva0iARWMTLWdvdn8Va2ciKlkCiSu2/BOYu8/gJ/ECOfNNb56aK7ZvBC6NOoRdGuXsomOQB1
6LkhM8Im0JE3dCZUivAnw52mkclmdPxCg5u9+LOaayGb0IkmlYQyxMipPfMV28z799rQ05FkeVYM
cLxzaqmC2hNOmXYeqogP2lW/fN6s5SRMDgCuShM968O9KVjs8FaBS3CiUVlilD8vOYgxbCvg87KS
brxHyuBltb8fJQjP+ArRCd5H/Y+1Sp7yrkgPfzMciaQFAtNUROdTKubNYFGIOnfft+MZUGcB0fEU
oz5eYmjV8b9jQulXD/fTUIffOgpdi1CvmPa/Xs214y8aT0YogAFRdmZo4G2xOahyadofsE9TvvFM
5pnQ2yshcqcjfA1LESxd1bFu2WKIgedFcsv3Z602q9My8gtOB2D46HqLB0SFfjykIcNYY9+TSL3D
6qPu4PEWz7B2vpipNSyokZZ+UUhEibO6CnhpL8FAbC9XfY9CDwBZ4v7aW3yH2msULGLjrwzcYQUx
zWNh332GtAsY5oRsHplskxa6CeFF7UAcOMFu+zJgVVDQHHIdB8vVnloliX/gIZ0hMYzK/uQURtAM
VMvO3ssIJqQaqtuGtWUPBCB/nAiYoaVvI5hWnCy7b2IZTOghDbiCRw2tc9mPaCrONOgFztQ8ks2z
88OsnYt+4kb3QFQcsmo0jLSXoipHFRFa7mydJiauSl0UATnD0pk9iR/mSXLJzN63YiZdfUDFYxsU
PwJM1/1o/VthhCkkszv1Ny1XgYoq8nrilHDYvx+3zhDHCREtktGR3aqf7X83RmfivT2hLq4IgRZx
d3aXHj320qkCc8mvBmqW0P4yaB2poKW1y/osyCaQkHl8u5YeO6E9zVZ5C9GjDo8diL2idlgRJNrK
eiI9LijIgPJSNlfzGf6cyrp8EY9I83G6M5lHCpjFDH+M3U89QKPNjzEur6jRYhlngh1732erxTJ+
FfDWCYujU9KkTlDD1x+EgEtjaDq4brVt/c0BbsvIMI+5nr9k2JcFPb6G9QMTEdsLu2fl5RXJMoTH
MekOKerF1gAULG6yohSTYs1muhCLQAXqdO95JvgQr1ODn9RVocfYPVjBsGzk3MYfBf1IXPR34QC0
j2KidBZpAL/YVX5tzukUYcixwRxDJjjvLsTDbLKrnAxRkNOWD2pVJEmVDSkonDUzzTFafzquJaAk
WUeBk7z3MIr73K4mI9+ZEle/HjRjXFPKbmD2XtsOby+w8V8JiT72ZzY+v2HGDh1FU7CemG6JHU8b
V9j1yVWqqYiUQd15V935KrXY5sLbGIPeMk9gkZxK7oP8VgAMf8QOa6V0hU80mG/KuPBSwsyHy/fw
lYqZrnTaR894JRC756Kbz+Xa76ko2u+n8aRKfiOviH5aypLmNd4Tt8LNWw6H4vKccNBMe4aGJcSR
WwAHS0pBv/nDz9MI0HopBcm3D9GK68Iq33R8LZ0Nw+LGs2TjRqiW3sAUp5TmmR1UM73CFkoGXyCO
EBmjxD2zBMVggEm8rbB/hvw2qJoNelA6mR3J4s6nmBlf1NbVEhmmInoPMrAMMlbqfBHXwL8uW6Rx
1N18jevYdlKDUhnrA/QmWxIF6wLIteXsN649R5AzF9sjqbqgocty0Xx5E3+Fj2QOkaxeDPNUGhj1
DgTtDjZWPK6EopY472jSsAqFszno6SNFnk50hIcbE4Cl+/vst6eloCpkkzuAziluxVkr9qAUmp25
0in4JgaOuRJUUDWrx3NuSta5Pb8d/ntAzkIiK5nj2Hmzc1uklYJoQFNzTHvQavK7Pt2Wnk64qP2z
drf4EcFPJOME0GDrESL2i4k27zfr/FJ5VRrfhe18WkCCXhEnxRYj19qW8ENFKclkfL125Y0bm7dd
GMna4SZI5CurkAPNceD41sJwZezwz58r2GSRX9WGXAonvtGq4dsFfOQZfGO3kl5LFaWBxFS7m4Bc
UHQ3/D+5fUZyWlCz8NKEgngYfXPfxGYSn6Kyi1OIT0myuuDxZZj0E/X+U8iJYQJZ1cmiZ/CBO8qz
T+81Q4UfVbY/gO2raBQ7439HaT/+zv/LyKxsSNWpuQ2e6wf05qH4BlvPcIfdvX8Pz2GUq6QIFdmJ
kFs+lb7YJFnwqhJcUqphuvTPGU1BKxXkY2zpLkocxdkFbeMVzPaBIAS98iUd5eAIPw07srqXePQO
mL60oXVvKc6+rpDF9dAIMaWsBwZ523t635Q6IL3HNz766I66qDXabzKsiWfHoaM4k3MPl0lHBVtQ
04Vd6+GfPf1zaGTVGBCgq9o8LXzz6Z3qksfs0iVs1jZ+hkBMXobA6sj7GyaO80tcZPKEO43eNHLS
NESiF3Dr+xQx6d10XbyfLo4sczhR25sdYRSgHEYYcyYy21ajeyTxxHhySFripRETJn6zaWl7rNzI
Mh56hxRp+3vfaq3awF6dnL7SduUANN8S0o3V8XM9SUV10XkoN+ExY4QzAXnqzjofs8RmS3mWyIlX
pT9sa283QeB6dlsIj/qEndCi3/q5YtE1RppScCqK+sJ+VH8RmkXwh6adCA696IefRmVch98QkVPS
JSCCOfUGNSTzODFGyIAf5/UdpZ/lh954tB1vOVuPXWZ4wPaQDuX8ocOEGifi7zSrqAJBzM75Oq8d
gMHnvi0J0o4G1HLGxt391jIH4lXSEMHEbarC+wRUyooj5CgH1eW8aaMPFHhHNzNkC2XytJQ0dHA7
4RxHrR4KHurXLMe//iFx9FsbW2GTptfhnXFNbgfn3ERQcox1c7NPPIu47+UGmRPTUC5LM0MzQlbA
0UlI1zAsh3KdgcwooqBNN6NqblYDpj5rN8CCutg1xmhodjL6ZreO9zsSrYMENopHoK5SN1MU+dYi
/n68SuP+WSv8w5Q9rNW8VxC/9SgmYxzzjAwOmtYOglCRcDUdQ15BeGr9F85AulsDYzegn1U9TkFz
VApuC8qairbAE+0UacjxYhcyaC/xUMOLqthkywSq0E/0MdshwIrDoGI3O/+CesMGDBccOcRJ3Gg0
hRIJzrgQ1laUagvECyNmJsoRn/GtBq8DMyBXLApF5tjJ74CrWvri66eqP9EudtpShXDHj74WEoFG
ILMQt8h4KjG4+uVoKyg3Sa9TOI5R2mOSEHpLSUSvp0af8pXJGmUATyRmXrDwz/iE454BFNooyRzm
MX+fAd7qSjxYfIuCUs+ANw3DZTTOWdDn0bnSrNV6IB4BEUeUPfy2c0kPU5sj0+3lXrLTAeDiANxD
EQDwaq1PA7GC+128oL5xqVp9jxXnddOpMV9gCx1p/Wf9Cg6b+JikTPQMqjgXLlGlVFsrUppO+eJ7
4RSm+WYXGKP/aU2meb7ny788fBLURA3rtJiF66iw14Wh0EFytSFfpZ33UZf6XBBIFpUxmYtLKBYU
iE/P1GZ7zKqftt5w9lNRVFsHuQELnXKUWq8vEcoyV4Q45827knbJFBNyeNbn5OLV0wFSYrEWfAP+
zrPBsZdgU9LSFsnNE1Dzol9zlflh1P8TIrRhjsHJWBDQdxg02ZJDsblAaLWrbPz7IhmitD9+G1zZ
YpAdmBUOf6WFCsvO0medgXi53dcz+WeomlhMgWTZq9eEZDrCtfq2HTszVKW5dW1qNY6OcUKHwe06
YMt/YyNstr9t/og+Y9zC2wAy5fKa9yh43EzqJy58EV8CACnq4N7AsNEcquy4S09j+cxG2CP3nRro
S1V72o8vuNV6ZMi/tiCOkEpBJeoKPO7Gg9EWuCTbE0FM9qlCFvQ5eW+h4HOGjwqOGc6jcJXDueQk
3ZebnF5Mt+Wb/0t+pzzz4dFTbufiUFiF2qvfjMoYynRM1ikf879m7lV7pNFFYwovLIVc2ysHiYW+
t7BzfrSakb7ntU/l1cHU03DZZCmnUuY8n43PH3ggezwc8B3QCTUT7heToOeIXRoaZ/R/UpJBFQvG
pADmY32Zj3WRroET6DxdfVsyAr9CxSo9F0r35HbI7p9VJ8yoMFR0djqHmFywwuyNQP5LlBXriBL2
XYXy3jw5G+T0qIh45EK9NyTUtHLM/GuRYFzFdnoyY7BybFW+tuOyHPKoY6rhmvJ3mxS1eTcznwnb
+5yrDAa6LLfJLiwmimnjb8ZHRH2WBsm3cm1BLoKS4mXsvn6IryJHd3pd9K+pRxdCUkAgJIJe8le+
g+/DHWdQlgdW20XogfMsSLJb1x7v7aAoKqUZCdugqrtmT5bRFp5KeiA8GQWf/5E1tedpPbaZYKTN
9Ir2RXkAc7/kjQ7r03PxDBYq7xIafOaVPnyH2Q+fmb5hiJcUyvN834i1ocKIIGkdRH9yfQ2YS2dj
V8m3W8A3QWcPKqqz/VHngXwtc7fNjDiqEg9OKnPwLjXTvBPg5FqHCQrwRg5JFYnWaQPnp8Gs2MnV
AkixRQTW48b6ebguxTS4xGMjSYSBkCqP0wCfc0aQDFm/7v0UbaOL7Brs+c0rz68FH/sVIWq+utVh
cXvtKkUUN+KdyNKKgdNHw1v9zOhsEojta2qZjnBo/e/X83XIcFxtGhd9NxRRE4avsJRGbA5Af5cp
gwTO6tp5pRTR0v1Uhiualr9054tNwWBkMQoFqZe3bn6LAKNcStfydu3qrhpbQbAL1X8JRBm5USc4
VfYIFQb8tlzoKK6SgCeBWRDaK1d2oWCA0O4t8PHvEYL0OUAd7bmfBL+1GYnNOwj8OvzVhwq4l/dT
75K8yR1UqJOS8Kf/07E1WwGKNMvQVQ+n3h3PEjlzAu3u5hUTxMOhRuHNaWZTtsyfXWa9l5fhVx1e
SaHYrUFMejFhvH7pJbAHb6azZd9JaaFAOGzjd5s4BlT+QRldY+T8aGWvtznKVYS4yXpQPl/WZVjt
urE751KziinROIEMmaPV8FJBI0KoBVeXi1l32l3iWKsfvPUEMNEo6dWsmqpMQUqOJ3KphKsp0L/l
K7l6s+NEEsl8yxD7BP1Yzg8hiSIaGY1Q4dWBzykARy0TALhse9Ms340wwVDtRp/jkceb93s2OXrK
8cxYOKl8BRhngwnOkvYGSUw84WHDOyQFQ+XuuzuxRwMqE7MdSrDeyxKQlEe3Anq4abL5ti9M29D4
wxoKLxAHkcAYruxFTv4/nKNc0BYWCA9MEgQAAUgDNi57E4SoBKjw//CZT/hxmGiTYh8EQDfVdTiI
LX68rwnkW3PY3cnf9Pnk4LM5FThJPvwL/5MXYr4dW/uTHaCVzuZMMdq1asahLAdIEH7WUC3SsZFQ
zUWA/N8YSX4yAWf4RTVthl3J1BXth1Dx4cDfdMhEE8ffmhpNeDdjNxSAFD8/0YTNt6bRnfZCwYin
NTBIYrweZX1XGVmRxOy2zU7Xb19meZxObFQB3kpAFloIFbYlune2HtVqB0htmP0ElwS8uCDxDYOT
+tAlY2BNXCQkCa2uBZOYsof3SQk4Q00rBuwF6dXRySsEUopFcEvbEkT2dZ7k+mOqM78Kn41Ewvja
hp71UHcgpBNempU1kFm0vSEHIDRx5XV9zVyiTeHNJFK1X4BgHaTK9zg8S2/CcPrjzdCAmsrMmUkc
PQjntx5umcK86LMlOalTuTeytBAJeBc08D/7Lgj/KywVP7IgUp2tPCj9ZlDvXedn2vAS5RPjbe7O
dyfCoZUnrGlM8AZegna+fr/zH3llwMrHkMfYq+TWdRvJeoRFANXzB0r7H21kGRdvWWOOlLCWlzuZ
be0ZpdGGi6E2lVe7dDbeO+QXhJewjcfT2Kln1y2ojSkxN7pYLLESlUC7w+2ooamMVIHCSAbxogLs
51DiISGphjZp+3iGERFwl5VpGJcs6jv19MDalOIWHw8BWZ3LE2GYyQnq6Z5wftoq/5/l89HiOPGz
UCrtDNyzHDvL7M79a8FDGxWyQIVvVtboFJ5ltMCXhPibMrosDAPdvxou+slzSWd/4ZbnSsIR15tc
JrJmPQ6WvQi4pDNVFIlyEKaXGdx2wPDCS5fauZfEYWyMAEf2zbsr7L5Cu0b9nUz5WiboXr0m3kZ8
xeTNx3ZrXp8j4+zd3yRp3AaRHRbmll4q/wJoPwyI6sjVh/ig6MJ4N5GKI8ZJ6jq3QBUXzaxNaPG8
fLjD8LaH78h1XIVxLYOqtV7helNk9YyfpzB7OjcT+8qo8c51XFSV3BZuhioqpsM8s7Ff9YlthFxR
3NJjAkFNnJFFwsWMw6sNB6t0SQUf9KWOCgZXrVYBJzB4eJRSa8fp+LrchGQ2eeIYgc317VYCISwR
hJdafu0fze6+9TE4T5Puz7+SWvoJuUDCp2UzRWsUJSoh7KMmXW0/XX6yPM9CatG7JHBWsGNtRBt/
I2YBqgGtvV+fMRBCsWmfCacW+1s8XM+BBUFuYFomHAY5GicOKN2uEsPJ91UIGUlMnC9RmJLdV1JM
ot6Xlgafu6sDqK3fQ5FPVksaP3rNNcU/1leQp2ow7qisxmcQxI35R9x5d7elLiYv1n5VA6wlh2Mj
KqJ9pb1D/DhaVojebjwGxkxTt/t7DxrSVMZgM1WKk5PCAytBeGPUwrlzcPosgr/o6pXJOJdD1I2R
MbUjhn7IOmwJ9S5me8xpGBVaJw/rFV3PnwgVpzpznXgHm3nL8IjUtsNb5WMGgIDO8YqB7RQ4miTv
LhT4SvyZTIFDw/0DLCDmmAsJMJAwYuWgZMrD2Sh5+suoxP+4yDgHZm65/w0acNmaH//vSz7/yQ3i
UWfhYW9I+WjC2c5wpTz1JxIYI2g0PY0hPxFVU7BRGBl38Kzb3Qy+JIdz74D7YMPuz/9IxQ3y9CBI
KWEuGogj9vZ/KCiqwwLjAbccA/FPK2VPz9KXWS3CXE55ur3mA9U3wNMR5/tZQqFDBZvlnuoKDk46
AfleIglFwQIhU3sOx+yDgaXR4XRZhZphx5qUagmc/3PNtEPTX2XSQSsZCWnzpu6leUeQp8isFgqV
5iL1GF8GIc8SxgMbzi5VfQCKRfCNT+7HLIjPlhmjGKJeCeUz0oXh35bpD9u2oMFjju+8Is75Z8kO
6GGcdmLAV7XvJF2in/Sc7evo2ldc33AQJkKa0YnJU3LTWVuqzz9Hd6+JZXVEOFIBbNRJbWuh4MD3
24pqWzypdVRsNvmo8LLsu+OLIkP7DN8Vn1TTya2D2oMJF1T38RjTOpUwe9XNpO0uXNAzKpQiKa0f
T4seCNsTGXCwaW243t6TREwhjM9KamqUgIDhZd7411HiuLE21CSy212c+/hLw3YcVWDZ/BoI4mmG
dQ9ts0UjWAWZFo2/U70KrhCgLVEe1SjtkUWXxCoT3chDIcV9YTSt0FMBfiFpTTCf4hYmlOTHyzhs
FxA5yiBc0uJnERwIcuFwN/7CVm/+6W7M7Ct0g4R0OdMtYSTOsXg0PtJPIAf69yS6vy/nUl6O4gCS
HCOSJENivblLhZCOH6Z6KixwjRNrF1TDSIHMgSXb+y49lrB7OGaEQGV9mCWehZ2JQAAbHIO5c9H6
Lgl6kseQtyhKiUUTrIzNVXir2+6zwsdxdzKyPyhC+1CUV0d9kNO9a10jdhd9aAbFQh1FPWzZE0Q0
/sjQifO3Qu2Guj6mPLSVUHcQm07fL9bVgQQUa0WX26t8S+6o6ZXVuWr3KCX8+M2VT+1XwLanxJFK
eLyn+atRN4saGXJ/oxiaKinTOBb/Lz5q4CQVhk9K7tJ8UyaPH3qW/y4EJOc0L+2OcKB2yKAR3roI
+Aaj0XtU4yYW5RKGNpM45YYsQLJXHgFHaUquUWPptiv5hFyZGPE86GLukx+L6f03OEJSfnrSIKuL
YgkmRSh9ezgsGWC3eZiPLUE8IlHIftxKt4m8+2I65hBhx9RMgRVQq6pApkzYPEYJxzLTX53ugUiS
fRm/PglWUi8Q8VbEmUb0WkHVwgPcqGMZfEg5Q/Zu19AvsT/QzqaM2377sEGmVxqK+caXbEEXBj2H
0Ulx7VsDZyj7MN3eQQpNjG24X9GzGWBFnCheuvaCuWmI/bH+U41jalVPH5PS6aov8BYchOlUjNT1
6ypRo+cIbR+yMDz6bmP1d+WMtlfkGRUJsRsJJw2wF6KPmf+DdbU+Vo1Y3T3MW6qnlLQzy6YIrLgl
b4Jjk1CJ0jfYj/Ag7eEGced2bx4xOCZyXwsVOMnFv1zPINaIHmHeLP1uZF5L+xwFOztuo2LO7GWe
z9nFjzkEcWM9SBSYopcab5GGvhxzxEt+cz0x82h5ve4cfRSQJdj8C6CtgFEiK1cIZoj5sCCJtUQY
2u8ByAy1Axg77Bw0v+f1a5qfFI71Vz3NKvxOPo0kp0x1T2Pegxxm6YeIxKzecLGlQ77U/htHGa+L
PMue20HXnLvTW1QUkEcNg40FTuZWQdu9oAA1h/tOLxnPa8Pn2uQkb2T6iWO773/dkphaQZfNBb9M
aoIFD10c1DQOmO5miiyLLovtiavmm1YWLV6saw7qb8ZfY54jvB6d5VrA+PBBej6fWLwJ9YTgf/11
R3SbXI8xvnTeLgvyS/TUn7dRGjmbLaNcfPbFVIxnTVmoak2caC9Q7mimz879rwU61m/gaj3W5hhX
EJjPUgImCbk/d66EpYtpIY0n2zAmGhlQU3q4YSrx2nlyYdSq6bPJrTLe/U2kMA45QTwFWdrwR8c7
mLnkoKwS9W4gJzhfeScb1X/GSWPbCDsliB3rbi0KlATB5gi4Bi/tD1wzn7guSt67gTUoX2kCvv8I
Y4c3Mv7VjxkxYx9/OFg/aoGMVQTWFnMDUMiD9rQCFPK2/9L6ASbJasqhZ2LkzPp5CEzO6hLRRJmh
pvQLy3ZRv7b1IWps4hiTL24COTji1JahL2x4Fh0A6/MLamCE+QVjvJ3oxRz2ihyyoaFDeC8fFIrd
dOCMXwSfGE0tIhakybbjy0pxXg0Fcgt/L+IFzvg/4QyEkRcR0IugL865N1U3NFclxopRIEOEWymq
tUnkUE4n+XCKyeycn6nYPe6rI+H1ZRaIzPwdBeeG+nJKKLnjmIfFC+wYhCzugPT1fTou2YD6eqp0
25O5z32EKjwCIkL3Mi4QYp8Bx9FEIZSwRaftGQR922l4gJ2jTDQklIFyRV9ZrzLn2sJghiWOv21C
k3GuMtzjy/c7QC3UM48UeN9Xn1Rv4FFQgrnUgXRxXf5Vg52iYBCOYktns1sS/LE8JQHUgjb9zgDu
sc3WrEKGml3NFLQJeAU5E+Fjei1H6PL9rK1N/MIEG+HL48nn6xM2h2UoQX7Aznv29/XPjKdGcD+O
yHFhl8hYhpQWdiZSiPo41Bh6p0F4CMduyRCo7s8Q11UyNNk6jtVb8ZZs9j1OO/CoC2ESKk71+O1O
HbzW/M2Uc4MGIq4EbF+0QzzjX/3hISOusU+GDX8wH2IISdF26NJRJPZPUn/i3wsNvfpYnOqa++hZ
N9MEK8rslMYpzrg6xp2VCMYXr3KIuSgeIZoEb8c4FBpQwPT/F4naC9+DGJbaxEBCgHSxJPjzt17E
pXDiyXta7TCgBOtUXSvrmbBPyS+pqSO7P2Li2I2xqa3ouewB68BqK5eVyAYQh272YJfE9iKU0z8x
hOx6Lxus2wKHd2GnEsAkNsdfdNTV2r8Cr1rSc3/OvAR3zNhfMvnd27s3yYpQtUgHJpWflK/QvCFx
uY5BNX2q+3jJmH73hcq21e8InWeUTmhFLiCxjteWWZ7Mz8bxgfAwIuVx+Ow5kvuJFN+/+7iQ2ZWw
/PJ2qm0HRJN4eLPsiOgoi/zHXerf6bXS28sqL6qyEwzYNLb0jTl4FCiaX2QLj8xHl+CNTze6f9V9
ECCKyV1oV5URuDEYrOtP6GliDw/k8TDv5JbgHlMKeZ7ti7nz+W/GAvQJnbesGhWtvz8etQQGUIFb
CfSruLiXREUxAW8hc5QOJdW0gdbsYukjiVm+o6P9r/UVEmOR3YOKQL4nXGLgowpoKucwBrZW+0rI
WmV430y2qQz29gevwnkwWKnkz+OHWbRjfs9D/P+hSutT6GXWpXs7MhAICKKwD9iSc8quxA1U/h2C
AXsW0naNUg8l9ZHmO8/TW8capE2UpsGfaqTr4v7Sovwxiez26pdVYX0a0RZ941/zv/v74P1x8zln
hyRrSTzWw8YE+gniFcMjvt7V4K9UA5/MO+pVLinyCTkPbt6DRrpZxT4oN3CuSXffMmCP11zccZbi
wShGG9v8wticizfcLSd8DGVb1HSF/FjiJTmXtsnloFf5d4x754ZFvK1F1ouxqGmxgDtT1e2AlZkr
b98Xd4PAcuz1PCxa+ZWGHXPWtTqSr6tAj7l7x4g5Lmgwuq1MSTsvLJgrdYhdgusI6GDYPh73rwnd
J8dh5w/nx/6OCBEWS6MN/tQMhju0eb7g/PkugZ7ADV28BpiHerfmfQ9Cjj0rQsPLGommLthrx2Bb
yKyPU8vqXc9HakOqwbssPhU7963RriAckgFdxxe198Ko9kJIoERnB4dMvyX1BGAsJaCVtsokLxtU
/6NsEyN08LVAH/yiHSc2BfVYT6Dg4dopBUDCLVhKSoqL9DWblkDAPwl1U/YeRWCEZWBRtpnNA0W/
5q3y98xmCANkoj8lZUXw6ht+LHtCKMem+89mQSocll9bSn6utgo7a/TXzx++LsMA8qQlkzLZG4QY
JOqH7sBXwaBueDRVdDoLCQkYS3nxOdfD+R6t3g6SVSvsiuk/AYgzuCN6GYUetn/EfENwmVn6qrxb
nQL04sRQuBzLghWIJlnxAWJfLBn44va1hjA7t+31J7Oi9mGcDwfgJ7KBCLeiRgq7BBIKXJGuoBwg
q7dapNVBnP/rVqgl6Ur37qec2Dxb7q2iCYFAnIL0/D2j1zFsmUMOM1fnLHwIsdGRbUrUTxCkiI/2
2mBO6iy1v+HNYutIct4i+Gw4LNVkI+tpaLNCdEXd+jxJ/dhxUAtXw5yf94zpcNIw5J2+oJQk/ENs
JK83IKL4qATOhW+MB+/Q3cNl+hbI1ZGcJz4SJ4V3BmIfhpN81cvvPQJATrklBU9Ltyavmhl6NF0R
2CG/+jZnNspK2jZ4n0rfZuudVq3cj1zZj35yxQ3zQu7ffx9gF4iLWoAnNZJRMc4ZF6KR4Es0r0lR
nzsjDuVxQCqqX8YDqkK1T04IkSCFLUY+NVm7I+0NBzYjn6cYSjKucahI2XTWw6jAY1GXJBTQP6wE
UHfWuEaOph1CWUQRCDz4rIbxe9ZcM6E+C0bAMF0cMd7DL0A0ZCrrk67qVcCqjkJqSgXbRztqAdtL
1sJXqi6x7kZEglCxj5kmxO2ctLCFocXQ7y5pOp45LS4y0da4V8rwy7UQD6yKq2iy/mH06+Bx3lQ5
I1nfvuxEQscfqNPlQa+ne/8vdXdRBLcCcC6w6XRA7nVe059E+DbqSscyazs1+1yaaeNs8eZd1phT
AcLYehzSm3nhgdYsYL7Aq/d8jY7xa0FXXNKrLJyrsBHWy8lJoDMXJTXadTCy8q1rLWPZt7IlW2tb
rK4DBSdEeoKPueVoCpYJVoiGdi6d9M+PdWr+706oe1IUqMG+Ane5FAnwAGdPUFHS8Nj/3uo5/q20
wwpW2FEa4/AB/5AZUZ12e8ZmixCBhg1OBpODqYK84HKkjbtdkJQuhLauuOymbqf1P1gcDqQZgfPe
SP3qxCR7m7e0a/YqtHKCpLqcAwiJrIsECa5t3Z/+wLUkjumfNZPo/+u7S87onGFaaEoyq7xwkFPh
WjvZ/ZEou/Ks5SWS6Vs4ctgypg9VLrBnpI3goKSLy5ghE2T0wsfXpDCbz1A9iilv5gtcnhECX5z2
uka3py+BSjTX9CatL2b1xGzEdG6z4dDlVmdTupuoWs3i2gywfoGpC6nkLSgDSbvF+d9Y3RgBfSvw
YJDJJID+kaXChcmOS1ZQ8pK447EOntsoxt2Q0WyXqJOfQZvVs3FvvTkjP+pRHJPIcyDcisNaEIqx
EK0yLaUuX+7Ze+iBG8LblqQrYo3jYztyn8NaNxbJbHJPkjuUNVymGbup/gcfM8pFM1sfxuX8YK1f
YhE/TgDAxX5xXHO21nFhrUYyM98SRaESs/eTlpSzg1riGslbOLcY1JmAKh/MAq4Y93KwfDUVSrET
3q8ENPNuBX2AqkUrI+u+tPAqS5jutUmkCQSbDjIhu14Ve6GEMNHWzP253YIGNbsd99OfFPDVZbet
HWQG2pBSIENGEv5HxJR0TF7SaoZ5chQnz8bBEFNM/zoouenB1otvgvHff2PwHJdBSdbOYDGGCTT8
GAEucO7b0qbEtnfWejeQbiwuDyw4zXDPmv3n/8qEwchmdBJYZirFtYai9hknsaYCo0iGMAHWiBiJ
0SYidTf91qV5y25JuR9K019A7dp4FpE/bgLD0l5F2QZk5X0kNhE5/5ZpRc3nQc6m/MwFk+SN7+JR
ubSpAhQpjeXv72pEfY7rApwoGQKYnQ+S1PSkbDe92FGWuED8hChurtyf25heH81xhe3uSUD00ZWT
PXPQh/2zhrtnZ5tDH8pVAIaCvRJ1802gy2HuRjykkvgba0WoH6fisiftln2K54cPYEIvOornSViC
6Mh/7u3tE0uTSqqXzlb6Wb+BvwJKMQfYqiaT8rKFzuhQ3NPMi5V/Tbw031knhKD2kRPVJJ02zWF8
slU5OF1u2sd27zEkVgiUu6V2pg74rZHa2LPot+gGfbyARlD/JaAhgTkgYfYL+HHhpB+Kx/aQkcrB
NAE5saRD50zr1NMpQiF2N9JZ8LgJRvcvuU5rP8A180FaqatkuR4Dg9CFvACthIVom4zYd2zzPMFF
kn5fXthl4Weux5JfXlibFDLWxXCalWT5LMBjoel1BgflvwGH9EBygpnjKPBeMY3oDkrZ52iJ+r0c
eecV2kd9uEyL9XxCwnvabldB5wY7s1tzjbIaVhWrE+gd5/58xAXQ00RdPY077TpnvLueqg1zl36e
60Sjv9OUz8AokuszbMF7APz1zyHageL/2IvzMnv4Ouczftb1MAqwBD9BnGW4zIOzAh01AwCKjmuH
wiDv4cCOWaAqpbQMMWgqm2urK4Peuet17ULFIzitQzJEWbUog29UOZgP2E1FSM7m9/wlAhEWU/Xw
gxiUx4MR3gFLbXdl38XzPrmsKyFM3Yi8cdEDkcFM2nY+eVdiyFUPlZiuOoQ9WcS69YFOywj7ZAyz
aVRNqU82+mUDtZM5u6OpflqreOyBDZGF1DoiHKSNPgaj6Hw5YEn6VUV4FmfiMp/i6KwXr6Htv3wU
IicdXuVz31cnzcuRTCe0lZWOojqpMhcowg/3RX/IDdfIeudmWHdOC6pGH7YGjYHi/9NBB3jGV2E0
9EwSub+p600ZMagfkSp3chvm2HbCQM9T1CBOOR85ZaUBkuhDq7Z+IS7HiQy4LOPvBfh3B8IfKQpb
Djzew0HqUilyDHtm6zC56NqWrqDL0C7epiXIQSjSIDpvYbAkMFeLuQIxjFe5Ap7twD2Bc9jFKASW
gSUqvL4MtmpQOl6ths8VE6VAhBZVU75yCnQcZ4/9Ni8p+EiCId2PyWHTZBZklqFvtkAMmmqls/Ye
IUoIQbXJcCCsDsYxGwgqC9LJKH8ci1XyEgm6pAZ6TBOUFnhfyK6K6qyx6Y1doAWpsQC7NtSzSlrO
7fSxG344StWgfBVcISILHJxtksVbkOK4m5V3DBplzdBDzKtN2OIb9DTYz9lWSspK2DVp4ewAI1/3
zeoCzoWUtFarlW6D+hvNQ5ZZ73zU5VpP/AZFL07GQrlUnfqFSZHisVbNrnQCbnOSSXcLadKqYbL5
IcP5al25+lwAZ90GvEZfJ4mdwG6+1kYLbhrUOmtziFtVpy3zYfNj2coA7CQUarlsGyomoY6gEQHq
pX20BG8EMJmW/uYbD6BKKygMZMX4Dyt+lN2bYO/x1/ztAsRsyxyTEuqCvzb2txVmscA1tgsBOqBu
lAibUVs3ws0Fv2dJ+mhQbxOjJstcShmb5r6TYpJZeam8iHc2YhQOTDt7bbio+kbquFjroomOFlcu
23HXfRqjmRRIWSRUxVvmDCQjuDgdZ9A7tSnjdisUeG4qe1VOUbJuCOjOxSoehrCyNm+JwnQP+8On
jkRvQ+RgzyzsNrBosGQwdxT/9I86npFG7TmP8a6/Blp7FDWRLZ6jK6YOU3ZVf5Zh+iQGol1Kwudb
KMXAb//Lu22J6Pp6tvQ7fjMiTTMoflHj2e8u9d4hAyy4opD/rUo3G4aCsV5XrFQ5FL3tiuB+MQIM
VSLjGnEEyJRX5i1hs6fTDCkHDyByz/VnLnA5BOTRkgT2RHB67kZyaXNit31CpCrZWb1CvqelHmMf
eNKC3r7+VOEwsgnY2/+OrjjDAKtZhnPfEOs3IfqQG2SidEMeE9mY1uTw61tZcn+XNMwGilTNgbbz
cx0LO87+Xkr1heUlxkRVEX+adXV9OTeWYNqvOahIFOJAuVGMgq7/ZrRbiqEHr0qOeSQp5NhFiDYX
a1FZIEQsizCdV8ChBADjFOLbsrArcidMb4Vda+2LLvOQx2zLSHCDoezxafmajH4wlMmS/hF3WkXt
T7NRdNNlgaRRQLrDNpa3uCZor4Pk3iADoGZvOnUREFDoeuQxKS70H7zUfCbtFt9+YlKEALwgvKdS
aIuEJ325nSkDDUN1nHfkQ9scKt1FAxJkkOKgZUUSrgtyrAFdeRy2t8jNTyHwqUG3+/qztAFjk8t6
5F8bN2OBuY6LRRa7zoNFbueFNLfGjdO6uR9Xs59Rvii2KExZi+XseWfLHTagwnFsy7QbTeIKuJ3L
XDsHX0rio2af3AjZj62zxoYmZupia1dGWJRWkcca8m+jPEigOOheEEleUxOU9q6R59AxzA8v9YAG
x0El3CXW1cTjiV8peQYgD7pOYYDbfyRreIW6/FjxxeiSIUmYic3Sn4KtQbSMAM/NA0dmVNCxOsi9
jNW1Hq4oyRIpr9erS0dL81SHlLQd+MwTMPZcYq477JCwWiGyj4K7r0WC1MtZ8iza+NRD1Ion66MF
K/9yfdIEqLdFjzm6TDQvtdwabXaxo55AqWg8vJj6AJ7/k+4jduuoj6ZEtUp93I1/aei3xfK/zucY
nxDjgHzIubtNHBdqD7PDALNb4eNcNS6DaaUJFy0fxJPsOUFYqY/9lOlKH+cBNEgkHvOXcFcF8zC5
ZFBFQv6QkMMLgYz3x7my5zxrKiMixJU2hgOCbYng3Zu5E0lxkYpQrJCoIb9eY/mrAjZFkl/nWSLN
9nd6ORHmmRfifoXZYEDKRQMB3x6sOPUzLvkXM7UiwEIf7pmKKYp7hA67MvLr7jq19r8cxxCcz9PN
ozp5y6dD0yp90RtNGmGaMSdAzos4LovjjsVeeVl3jdWW9OGGihN2wNCe+enOKxPVzTzyqmxNiSu4
oako6hrPlY143iHx9iBl7QlB2G6rmiTl9WJ1xg4piDxtTMgCrBDb4QaOPI9DdbZSyZwB2cgP3XGZ
dgiy6YmCFtqLfMYOczLP4w3IRwCWQ/JAxugY/S+hkWr21Ea1p0CG+9So1FbVVaGStEMZAzi6N5Q4
0P8IsWgShzDIRC1vS8YrzfeCIzDX9q3n0zzqs81JuJ6ioqL5wITXagKcTxIGFpADZTxcljmiGpm1
NGB/2CCI+opUd4VG6FYE0z9fOgsbyAMupmECNCiJnF1hqi2ZRKsSNfruU+jtptr1EdbvpeDbO3LI
ghqBG3Eqcib25oguvV1ovrlBe59GXyc2xUZSjRFbrvxgkAgkMAMCMMRef7oz8UgnEf6XPrFBMzAL
pcstuokY3cffUh87HH579t2AjVVLUrcZZFPaG/CBCcMWmMjSj26DXqr3pzumQ87bXZXtpnLe6HNu
qoYs7Y+gTmcRlWGZRVvbPsFSXmLGXLjqR4lv8/DEc8+QFHfEN8znqhIVZeNMbFSdYEXeId3tfFrU
qUT70aq8mxeyISzGDbE5gbuOLBj44E28pPOXsZIvHVvUjJrMMLTVwE0ctjtdcs18/2jugATMbJWB
muG+WvuEOC3fHuXKIZl0ARFUYJT+Hw8L0+9rYUe+ZALtY6vZQojUtjtPq5NZbh3NHA/GTJ4BXQ2c
FwxwmIOIz5J9Pwg9449iN3NpNC76K6dLH8PIA/Et3CvxAQFFw1OZOpVoYyr4QCOd2DhQXhnsN8Ei
cxQmYCv+yy1WBbGX1SJURWY0wrI1ESbYVTUNx8LiDqYHgjIR7t05mXQ7khcEEbw4+S6an9yGfRgh
+J5eS+X9l+LruBqoAopFlB4LOinr8alx+bo87lH7FSm77VgNRWGQIfq4JdxAuD8g0+MkweOba/PD
4jYeHohXRYQPXh2vpEz+OhfXVxD4ZWp+AcE2y6vl9Qch/qlkoU6OXkj4Y/j5zVXL+t45PVyF/Onl
3mg0qplcv9Uz/x0ECGWyb5EESeueFesvOiw1SjsNeZgS5wodJfyccqPJI4oWpl8ipAMAHmYMEYHm
IVOLxwsgtJ8NO1iz5C6VZ1vKaZCRWeJdIlBXVRzj5cztHEixi8oBDXwzWfR9ov3+KW3b0VjAB60t
Wbm89a/wuQvu25q0tNPKe3FkFpi5tlVH4IkUHeAzT9hDkP8DAfN26+uOBygpSfswcpxIvfVXWC1n
gXOpSx+bIm1pd3NppIGmvTsUjPKgF8O39jsXm9i2TokVtsq1SujRnTdPVpSbk7xcu+ar7wTaJhDJ
lPS8PpGdQ+SID85nDGVPw70FGmaX3PEdxI6ZxkMt/lJArxDLZt+21K0kKj4azH0VKaeuIReQeStV
jib0cTY9nffcIQ1IEahtxpsNa6krGMYtZc4A2YApHU3qDC47bfeLOJFmpRXY56yr10TLxlpZhF/x
yMMQwtpniwf+/ZS/l8QFk8UB5Inx/H6lGsRwZvqZYVyLH0WpD4X1Dtmm+aiAT0kQCFw8FzhQKkd4
CO9zle2FbYhKdx+5VAapa8nXG7POHLStZwzgaX4c5j+pKygDFlH0pdwrlZmS9Qh0GMS7fqqC1A03
nGJnM42tyuxtKzM6tp4xVRYigiK0uKb2dqFYB8U0cSoYKbPbn10WqxTtJE6QglzwBQUmzqb+oIiC
Ew79F7MLJBgZDhX2fG7o4mRECCA5KFPTONrjaYusNs/W0aBu/U8W64XvaiyGzzYSj1AcDjua5zZv
I38p2VvVLr+vd/Jr4/7REF9dMThStHKbEmzjop4fV1CJZqHGXiSEsB+lFBh4fvufwcDaWgpaMWsY
aLzNsjmED+X57ue1scrEAxmJH5LQnANqeuRpLFKN66b4XPddngNBJyfyUwAQNgRosbbZ+yRT3z00
oamtt6m/CaW/M7ADl2cjJpXQsVz/Gt11/GglMfgicsbzENpfxg3GN/dmFwXUpbYcR66cAecG8KCf
+z5EZ7a/i+mT7RMOOOo1WyxeGXBFr/luDYkutemelx0yNckyxdjmu3dGIlVuO5gepWGjliz648av
ow7oU5hrafu3Lj7udTlTNMWd8zJme6/Iyh3iXNvR4fJ7+YCs8iiZeTTFXMEppMxak6deQIfeA6kY
F87cKclya6L+eXSjsTdvLhqIZqGCumBqi/lWPEq9zu0mPXKmRq6xPfgc2AUsC0o/tnyWvuRXjsjm
2tnGMPNxEj5KlZKuljOJCHswDr+ykaX3MilaS0+qMV4ybNq8ghO1xDag3X8AS2LmWtYZaeOjI5yx
6LrFAUfDwJbHy8wJDhn7zbPCQ36uWXiOYA7n82YXlGjMKhTIPaEqUaXee9cCdiTAZRBM3KY81GQF
VAzWOLQMmb/FKbJhueRr9pRwwMpnTSkg8PWe87A18mtRHE+Q++ineqqNa5fTm5C/61Dw3mnsqcBp
RwWvHHIGPP2c5jcnie5jFMmwVgp+nMidR09ty8UQp1rQW+QdF8ceB8LyTFPnvPoXpEQpKqRJKiqC
HE1znVWPIr3ivXfqczYosSF5BtTsZRgsSq0k53PQgdgNd84GYjS7AjvmQJUJ7pgdsjsGiorvMxUj
2GN49CMBEuMy3vRs6sS9S4mX7kVjAW4YG+Og161SQsZK2NMR9bdFFXtu2irhmlf6VADLjllZTxDT
/M086fN3NwQBp2vZylZ4ywg2UB8IarzGPJ+93ssQ0VDEsNsEnuKgyH/llPdlKKeUz7URkJfVu++G
X2o+9jVTzjY5Tk2R5pCrVUIqltXzU9NKnHes1jTBJOCc/SFp871Zny6tZgG0EN993m5PTLhCua2P
fJxNoYFLHFwNkUkmsIRV37wh0aR/bPs6e7o2DabGaMDQfM4hyETmxvR6bm1ZY0QhfPlujRmJochC
IR2MgsDXVBgY6toXGZpg3HmTnGZ25hZPAOCXNBmxanhfccmo40NQnIGC2sG8RzaPwPTax9Ro9YO5
VXkO/Qva0Q5aQdqP6/ZjYDXgulsHiz77StdYLBnu8y/EJQ8G4MaWi+N2QXL2J6ENPNihddRQD5jt
Xj4Nan+DCWCdQKGlncGiDpg326bon/4ZdV0G8YCY68lsz8mTNyMx26uRmw+5kibdd1pMG2sgfvUS
NCBbJAdTInq/I946LsZ4ak3kbqEEXg5nKktRXrAdftdT2CE5cEEemKQoK8VFbnnvqpYCuSqh/lci
shoc+tUsBfcQ57QYGdrJ94EYjxdhCeBvbkF5FDzkTFoOGj/dieqe0kLXNoK67C9ej6Bno0g2eGLJ
OeRg2NT4SILtTS32e0b4cxgnetsGS6kIEEIzQNoW1XBCfvtEs8n/lKdOlqVTDv+vmS561uvG4RQG
mAAZyghBYKCpDNz8LVT8mSAYU+ZYpnpb8n1I9doXVPsxKkBYawXHl857csm1O/S7wWPkpFPhJLMS
FatX/D523eprtIfT+l+f0x7WLfION0SdQGdoBNrErztpCJyRbRzxYLV8007v0BZaHVCltuUQav0V
nOfmMdC2gxzO1X+sELJy5UDQDgB1jCT1sp3OoJhltW+38jxBWv8yzhy1EImRg/XOlUy4kLhPEUTI
nu9eom5bCnsVr1KMACJzwg7rXdYkUYIgi98gI3M/d854se5XZFeg0qF1Y9NdJczT2wbyJDAiE52N
x44V+BQnXLaSrqgwdmbOL5TKG0vcFzXbqgYT/JAcXlQOIzuAScoHROahwVSD9ADcHIN3cU0ZpFs4
XZMQm+NnHUjFtuOx21shjzqItnE2LWwkK0MvSYUAmFhwd1GnCA51h/6fqaYeJh2cLCMTMnvwjdhw
87agDramOpFFhKyLVnUxMczeu8a21ACj0rwWR1vJ/gz9FuJtMrFLllcXspWU4MFlKzmta/i/Kw0F
MOsvxvV3F++GOpabs5gNEdvjTgD0tXXBGxXVVqY7dWJ2mQAs1DS3IBVovYKr8DyBK6TqrYfGx0wx
4EPk3wn6GRJ8U4gAEjK9JQ8w3Y963IJPuiJ83W6g5Qkasr8YECVDYfiJuY/0xpN5jzmZ8eRMEfc4
cfCKKcjq385WgCJorhSYizxPKgMmVkxrqsa1aUtG+j72XLDKM6BxLbMQj0sK6fUrUtSVr0MG6XEB
9bJvXOL/RLlCbYZw7NKa/FIPCoe8QXMdKE4rukYRnFS/tTQeqo93+TPonfTZhtG1o++hzt4K1CY1
W3at8tq2RDjcV+GoOeqlIFJWXu9FH26NQIQBb/Zf49mlJhLujGvYsyPKU+mnBmEn2xKD4+GvdXdd
5onqGZCP7Mlfhxw5YlcQ3KFveZG+DVnZKKfoh7CVMl0f9v4huLSvz06eoycSIhW79Mur9sbTIU2L
OGaPbzl3oav2U4j0aAEwzElvdh0PQtLksITxp59LYqdZjtmqsgHLl1xdvJ5hplEFRNRso/LUTEF5
pJlBzCOjMtlYptYLuYxM7hAxk6aL3v5YPeF96di9GnzdEQDVQUU5v2R9g+YYLdp5cazN8bFQlV0j
sdiKalQx9gG41d4hRAQWkaKfBMiPziVfi96xEeSMIK3AqohxXOpVuIZl9irW49+nujBOQATDscqx
1DEeTxO4WXesIMQexxxKyF6u29QfT58dJTyHpqjv2uTf1ZF6PVHDZOAVjcJOQy1UtIGuKuNZX7+T
gMpAb8Gm0UNWpq3vuMI5SdBhwjAu/DL/Pf/Dzj6JjWe5s9dOD45g9pFXT/7lcFKsnVFlBkZAtO1C
R9WsCn6JFxNM/MNxb5fMKr2e+kNIK7vdNLLTfHPkAYrv7qiIpe1hBU9SHaZd5lkmZ4kyCPJMw+UK
T/0hLeyHQY3p1WI32BLlg4NWf2tfUjiIGR4PAevkxyQvjygc4xo4CLn9ViWwx3WndW9CUyyFlH+b
HTtHTFRubpmKVGsoKXnmkspZ20vpMqGsspF3qlafj8BSJP3h9xyAE8MJ7PSuJ++SX1ixJMJLvaoU
9xqpVTNXBbP5jEaNgQPIFUVZrEV1Xzfa1LyJdQDRwX7csDbz8k8a3Wifw9AO4dDhREq8Y5MbZJp1
CmARiYliF7WXXX8V0IUO+jKnpK7xb0hskOlJ1pTnqm3Kha0zCN8PS9vv0cio2xSphv2zNzhrkLzu
P26ny+KmMEcpVsc3GwZS0CMDyQ9hF6QdNDYF6jgKrYQUZstQYKP2wnYu6Iimz4REwPifmRR9DN7E
7GEVF6pX056WPA5otj0M8nTsBaOLn6wMDDGvcfwCE8h6zxj1RhrnY1pbr/WXa1HusiFiK9bjYBeb
ns6ceskn1cEWaCclOKm7xAvo/icFj1rbGFq0cmW5FhRodRbwBR6/GsATcA/bqF79EsoikK2Xy3CJ
rDwOZkmBxGqUqfVZwtwstkTfBGX8J/5JTMLyJmpIu1/EP2ISy8HyJ4JGis6l2DBzmuWG+MXVLkfg
VJt3ftUHfJFRhDX29clr6VTVqVJ59tc7pzzADqIUswkbl1Wk6hqyYtJYDg9w47e91VIgeIKcV/ac
0Oc/1xm8aYErmJ4frUyCNNIqqn1ZF7GE+Z3hqFUESpfYxJqbFYmfkgPOadFVnVs1m7MkIAmSeGvV
sfVolEXKqPjBASlhnWtEoJHVI06Pl7bV++fSSuODvVgZlLULqqIoFG0FRTjyfRk0gEKClFS58ui6
9U3gd8rPGCMWIWNh/IVcViFbq7Q6Dwa/6Mkzu0PtI2+Gd0lstsViNilD/2lK0wJUUv7guhue6YP1
1LMKWK2xMgqsIkQY8l3rtIg9WIFB4in2In2RnG/8xw3ZU9JUqdvEflkJhTlXqPBK7NJhson54nJX
rHNxwFfrvNb1wyB5bn49CK/gY6Y9mMyGMtdnKL5YgGd5vdGYSEx7u24tWcqIS6ugHl6vA2kmV30P
loHVabeK8vIJpSlgHzru366/VC52794pKEehUyRns8NLkZwrON7df8fqUHSdMjXhlF1gQxSAKdN4
kpmi6kuuhmDzWhzwhOyrok6r3e/+BeGfDz1iBTITPIoMLnmCVSQINhaA3q5zQg1Zl357B0i5H4wD
KZOtW4wKgNLh/4eW+IbN6ukWMCTQgQE/nPWK/83y+zbU9EKECz2UShNfW03jrkgngfBzAEEVgE8z
xAo0b9Q8XE616W10pxJUcVgE0vYM9a+44cZuREzn1sLND/9nUsyW+mriDVg374bY0RWKhPegYDAv
GdrlTnkSwkNEUoK7MknRssFggpqRsbZpiYnIU06uZqhg0rTsxe1M+Pe7bY+cDJo/WPfM2i/NMeVe
aej5HLTFwkiyQ6L+ekbEhwdry9Xn24eg6GK/ZlNonJ5r+SOiiigAonHXbiUEF5BMdK9xwjT4zkL9
3rC5ApUmsMd5OIRUDCF3sjMiz6IjyEZXhE9cTpLP/f2NePbBVIDhbVE6c19MhoDuzrv+Xn1xMmDz
5qBsdeEgkW/lCtYtqQexFxe4lGmoay/b8raqqHWyUjVBgsjsRcNOgZcAPf5DhN4X/i+9GUcLMP1L
+Z/MonNhUFdEAHNnB+P/GGTzmy5CQKFeoMb+1Kpu8GglHpmBk6YHrPjkBG4MOWZot08oZnxpVhsf
ZPigLymz1Fv1ThMGmnbAO7hGS0f9LJru/eRREutc92RJE90vZFysN2cu/Gqrxj8vos7hXmFElRXj
niJUqKh8wexU1LnnjvqwdV5YJJ9xjXkdd2rO11f1ChOCFUMwD1vWFHa0D6We1ILs9oAS8VDAa16J
3Oi6JkV+lJBqNwaJ88vKm7VC2mutssX0piBxyU4N5ZOI7TSEFYdSnbAfNnC21jFWYRexqvFrp7rJ
brNUcd3dwUzlXK/m5DWKNTEC5KinahnM/QdwQicpWaYMkXQgRDNE12MrMsgQLALEHt4LkfR78dt0
d1U7BGNWS9p0HtE5PuL7M4KJPUpWxSIIkySQUiDV2UI6S2cdvPyh9qbYwwqs6R5LUcAdaf7EXny5
sCnnJ2bIps07ufm8na1N8vbHif8I1rIX6iv5E4iq370jMOR0j9p5DZNz0awsG0dgj9jRqugvQVTB
7IfggucZ7ldz34JRXFJyn8xXLI/J/GR8pUNLXulYHytta+yDcPsCp/DzEIHQRvK9Okr2a/87LQ06
MTyHbDmm8jVbOdIb1LnNbzp5vmAgnKL7b9y2iJX2Lqq8cWh8XiFj/eoaT10A1tcTHEU3sMYQy1X6
2R6oojDfmtQ4cx/akYxMAIGwPcHILgYTsrevS3ro7hWkCsw7QnV1YKeQFdLgB8gQkF1FGeYUPj31
keuYoBg4rgfVFYgUtLCzejMCGqXzoYGHEl+Vaf7IYBjX3tG3BIV6Kc/e7dkhpW3ujqRHkr5RuhRu
VJ/6jpX7iUfAyjJwCA0aNZGq6YhlBX6CvsSGYWwEuXLERLFQchQ9MqcYrHoZVufTLYoTQjMDu+h8
c1CTRuCLqQNBCiaOE/LsUN8SETHEhJfL6ZJDKVoAo/+ha4ljbb2cvE/rgXMmqIsFTPduFh8PuWBX
y/v4v63H//3tN/QgQIq+hGS2b8WfRUjjQ+Okgi+dFLDRSawWrEyzdD0et/5jZ8L4G11h7nM2BJdC
THcf8zEMiWCInEypB6xSlMKkcEXNWSQEsAhg0+kU+2h4GG6vXyAwvHjmBQ/CafGpmulLRUXmgshX
VabS3+socK627gRq614zIMyTKW6yK8KDVg9cjHWU/zfyd2Q9wSGSwnTAFc9DqdelSrLfBMce8x4Y
JKn7td8sktJ+dCeSr4Zwm8wiEH/6iZmuSEGuXD2C+18Aw4BU28NqD/cYHsfU6CbgVs5KzPP2da8v
h3ckeaWxnuX74x8Q9o8fo83f8VujCIlxW1b/zJrR7y5xsnvr2UVj/WfoTHxQzZz2jshWYDXcKNDB
U7kiqoIitgqWC/KxE911N1O9318aiDxq1Bmzul8b2qMSUlxOwc+cuofNx2MgJtiWjGSeYyfF66MW
hiSntGkeyJMfD2Iod5nf58y50IQNECcOo9aKUsDLhOZeJnTig+xE99ZE2kt31+hoLyCBzdmmf+v0
L8SZENMwuUfLBfkNKj0ZQHBjJFT/r9T0Ac3fC5TVdOW+r4T63etm4KkiplCqhakhgDPHVNlkgluO
0nkKEX0jQf5zp3bFNHxnXbCMifMNdrVgZeQLp6T1Vrbf9qRv7ho+eUn664iDWN4+X+DeAgqbbTv5
Bqsttr9nayNmKFCH7c3E/WWe1g9QFEAwnZyfqqNCtgVrP1lPmCbUkrfJrGabsol7c2tAFhuzHdyM
535+GcBt4fbbfrdq29BkNRLZAtlDKTiHSlubqFBu7LvNb70eWLAwtjseLfgjq7KdumpLuZxWCkWO
yQrss5OJgWRmzSw5AhegAurCfCpmkFzGzBfGduEeZp8ciDos6dc0nIf45um71f+DCLpGA33Q/um6
n+23hsKJ9X5b7Sm085s93r3nZ9NgzSB7mE+Xx79UgEStKgRuKqk+48eJpkJ5ipQ9SexN51CNqHqw
xWDDBIKCUYg9ad5/w5LEwQz8veYgvon3CaoXFS72L46WviynNfhr25BYuQupOeahcEnn9YsfKh6X
JMF3Y0Qz0YNgUTU+vdOq4jKrcrjKM5mxKpCJA8xV6sBhu89sTPXNel6B9AsrGdc1/bFyiWRtzFdX
RTKgILrcR3lQ7A2My4h2jxLKp2PR+esPwn0KZBAgbFbuMp8vnnlIcQ8o4r4TQUGCh9IgAOBtAiV2
vLSvYNpA4jcg7fRr56U4bUcovTouKZIf2i/jOj4Dp7jByPnboQC2BtsNC84kgNnCv/PqXoDfuFow
Zezlt++pDFixoLU7p9riv2m13/Pri50IdsKoumj5G2Vujof1p/ddQwov9PwvrudTm5P00ij/0VT8
kDz9oiyhNN+ZI2PclCPGQB8mmbxMhayzwabZ1S3OOm3aHLNwz7spk0+VPXi0VMNDuNJ4Vxu/Jjun
Mi/v0GsThyXAW48kvcvnJY+eUQnpLCWVkXk/dMer0mc5o9Ay3XPDTBvDnRvvrqnCbqCyDE/4D3mE
fX0RuJxKeW6c7wV+i8OUvrWoLW2ue9SDuW07oaTCRqJbslaf6UsTeuoRFiF6QipkZXBS2yOJdVs4
4DAMYQQXuz5fvvT298UFPZpQ8gAlScNB9jiI9p2p/VD6Dc7mroD/7J483pqXfb6Ya85rCvQlDJCc
xvueMwciRIfjV4ijKq/uel574gJFnzu60gwW1msbLql1mxvd9MrXHgaqiR9XDJBJCmmEt5TpBowl
rjQYYMHTDN/Z4vdG0ZvWL2p/8+JsbvrL5Y8H2zgklvBrg7pbYovNlYbeeoA9reb6a2Sv7rrEbZ8+
F9yoiA5/MtqOrpPWG/Mh6R/0dlUvH2JTfWJwpByTY4Cu9qsXc/DRYjHj2ucgU3IuiRZGH380SJ6y
0DLN+ac5q9FJtOQaiWNII+XExgn3RccO6P5Il9hwtwEa8Rgw7BmgRcIcgOjwA+aORwrjPrV4lQZz
xHm5LfHPqnYWhTTrF8SO9E/DHMjXgCNv1zPWAWay20XwW0TQkTrwlmpJcmQ0D424/rZe+R1kPb0f
MKsed6wUPc8hmGix7cOojADjnhkgfexNs2OQPF6trGJ0PGvtM3ykNxdr7CpFZoM9SqhAdvl9rsd3
yk7X9zOVKQRDrU7na5NNsnVaWFkmSEGsGetcmfVhnNhGlSVsc1kIPK9ufo2GnkCEgmQWYh8aHGB/
P9qHya9NyiSQrqCHUxRDWH7nYUCAvu4dl/k5TDi08VEJ8qefyfYxo3Ztj8ILrcB1LPNox3PndhnU
yeT7hxg9nky84HAmxuA+6FfN82DvIl36x7M4xkCj1lFK9cvVwzVknjkB3ifx6vogXfG2/NfNEPkT
uKM8OAVvA+Q5MyMc5bNyyF9IavMfscpMeCFSD5BXHUJWN+P/TdJ/mBP5BC8oxdFM5iKE6RHHC3ms
rToYTnny1BhHFoKkAMN21UKgT2Ytx6PQMgckLZFIBKvcfh+rax1ewBXp5/CnEprR/83lQjZWYPj8
aL6huRj3364uAV+kiFu7tMoLK0NjW8Pcuy1yMzRahIpBKmKYuZP11Psv7ImHnT788BdwR4DAJWsG
hWuB1B4r574ogiPcS9imckPd9TDPgjECReTM4scpyBReCU0sznZ2FSkAcS28XtTgAs9QZCITNI/K
wHOoYYapJc7BrAM3fNKLI4i8ggSgrxAbfSrw6U3xDn7MVkg+wzsfWhda0itL/uufD0uhxLsOYqRS
dWjhj6Oy+4VTh2m3MeGtOpT6gLq33xy3rs0xmxIKU3JSGlj92jO/VgrEuuTMTh0MkWLQCKNYIdq6
unu6MA1qldxKvhIu2mNdE7QqO39ID3VYBVjrRpXnpRcT4Kt8g60ytbRlfpGvB/cF75LJyBjwrKtS
ycasRXU6nGD0B4zhFsvWsMcx0v15vA9dG+sYHm+y/p1JDUKcDXMmOzb4eMBagvgougNwMCwUC5aV
eJU/RAt9v4E/OMWx6LVKsmHSUhwkAQ8SbXgjmJ5/ZPL8RBdYO3lCPJm+/u/8x54Wpyg6dERjV+6x
GrIfZQvTPZ3r3nZLSL+0OD9dsbsPot4GJcDCRTpoVoMgWMelEXU4amhASFoWGby1TWAem5xgpdx8
Rs6wySMyf7DSGgCmGxCvwTxKq1WPB6xTSuS0L9QsksH/SC8JIyxjFaLWM/THdGEDQ9qd0nQJXuCh
ha9h74cYSuSOs/KoJWNpjRRUNXlxnJfoycjqMkgdehVA4DpJIA6J05H8I3uBSbxgWJg5z+7HlvLB
uBoIn9EhDRhDaK730cqkUfNe1oob4n5K4gWmZuj4T9kOvfcmF9tZiw7+71wlRiRQj5F2WowfhEG7
Paw4bk47JZ0tItFF1ucG8+Gq54oNrYeFiT95+oeMQBHEP1jsaFAI8JLoPhq8+Mt7CrXhOQ23P/Pz
GUepC3ytw51NHDdhzOuojsPrhyxI+JhGVxtFVfV6P0K8N3l4IRbybZugmo0OPwal9aE+gYzYr0uy
gcXh2kolqK2Q/4uAe0Kp3HeDDXPzYgs62NZZ6Ecx1roFRRi8xaCVxb4qTMzN2kD4ulKNwh41OT7f
VFRnEJxTNLVm/vIs8CEg5fwWsLoJ9K+As2iFJl8xeJqS9HuMC2WcnjrOSYHZ6yfziiHMj+N5hdw4
Tddd0xhOPgDOx3PQlOnz5MShcPfR6IX27pLoksZtEF7KtrmiPkf7yRwivL768/iXZZg1DtKbb1lA
jsWkeLY6TtiKppeVPsjWcxBntDozHKLf6jiEVLxYJyU4d4AEU7tITFUKBdUdykv6Rb3INS1ra1BD
RbXCTKZesLQJuE8uoakg710iocvlqfYBWFeMsi8kjyOHm3O95mh3TAj/sSoo0s3kpDfDVWeTyjut
fEFuY6tLVAqYrnVO4Wj1YEWNbDeKXJckR1yUdM4zY3HJuhTjI+WtXKHYa7I3+hHncoReX4mnT7kB
laVeQNM99z48U/43BLfZB6xs6jHFw6b58wT3mU7o74+NItCOIjEHVWbH2D9ViCVTfI8VThTNlmeO
qp6wdsqQpWWchv1BPslO43cOlnqbkGw0MH6U3Vdn4YDSY2Ot+w0UA+NWVVXgbsinjI6DZflbaSAS
iMim8wgd9qnHRABSXK/ZUiIMcYAKdFhMFy8t1+drPz10fpaEYBTsa1DKv7cE/3dOIsSdr8SLj+4c
Yu6NFPRCNYTpq+TVMCz/bQTq43bf2z9KbKKqNzAsQYs6lFdE8VyQ5ydygcQLgA6dDwtc2lTUso3K
0Abm3DahNpccivfTRirKuaBoO0zi9XI2ZL3MBOaOnNvIz5vXxB3hdKw8IkuuCmnl3T97070Chm4W
lyj9tp+cJe55Ty1YtUiJNrvKzIAyvmYDaZdR0VbCDFZVqSFLd3GvolTxSVe1dYrI+3vqvGqL1W5B
ETVXCfoNrehyzdOtyqht8btv4zzuiktlJPyh0UNS2DtTMCO3RcR1Nx0qDZc8hatqNv2oWfj3kAk8
Ag38XJAj4+/WLzl7j6P0i9tJ7t7dIJf+ZZdJSDp/xqYZJVMf49bTWt00PzEbLyETtJZabgeVIAtl
fqgJOGxGXQRDTkdg7vX0ibH4tLRjv15UbTlHyCporH1kj1YQdgPIkfrpVxkA8hXmheMry46II/6L
J6si3RQtyAtZU8fapCCJb15bm2t6MCWXTxSHHGdEqj8320Y1GB+I7a7fRkjVVWjVcV/pYAcKuvn6
Cx1k9+je91ywAdgBmv/7f2rZq86cO207Lqop8lt1Q7+y/TknlQAtUTvJ3Hw55hu3qyplJfSIC1Gx
0++ybi0/aUTOV3DNQiSf2+q6Gk9A9YPgEPR3kwDNg0gRzptUI4CNHjdck/P3AxkTpJKioN9tnzmz
lqKz1FjR/A24ibBzi5t8uHI2LnfSRkb6+s4lDXSjKeUpLXXsZFNe1oU1kmW8b4eckes3aC8bf8F8
8229toaQz/Pt++bgn4s4uWCY1zLlCq7li4A7wZ4E9kUVZZNHitqBqXWoJZnBBXpDUSEnojVyvleN
bNx5+52qy6Dj2JA/X13WI6R7YvXlzwOdNXhKyXT7Knjb2cmijai2aoukjV+GY++Xvl0pWZd4UW5J
u8wV/Uvhj3SaB+g98ASjLwPF8neWzLDWRwupGjxLXnl+sXnqzACfDka3IUjY08IhwVQQeD3Sq+eF
+WCbdFNU/WNNoAJZhNakR/sMZfNe7iK4CeMPA0h0J9gNRW028IjEYnnf3/ERcLlYoOp9+XUUVXEz
yQpLpxdpvMKXK3SIiZ5ZVZoZE+MkmOdyZCckabnTVhyC/8LZP+ehUXU7ICm8ZHHluGixOT6z14hp
E8gjR34RVvk29QEOCdch15s0cLLwKClMLN0fEmUbUTTt+Fr4hiwfkejVJhto5/8CLQaEvjp7C/wm
EFNWYxWLLri2GgxraM2GBXnRKCd6Z+Zm2kJl0PVlVYhvfCxdncKNlzL7xBQU+tFmUXb2UBXQbDB/
7TvA6XPFDOl6eZVCFUDbsjFDODIbQLuNxswtH8j+i+w41cymWxy2FEF7nUdPoFxMLzLrb83wwbcJ
/6emw+bKSuxx8BxgORNjGdA2qKi/3cg/YRpIjjE1ncwaxWQQbbQ/GDkDANhv9HkuZabGdFebolzh
aYLRKJ6GjY6WSwJL2YU+OBzw3Ab1ZUD8DLFLA+A/rPpNiyMDTUhIQ7FFrJ0zU3wB+kORUXKC5Jen
owEMV56K/hI+YKoGtPMsLyeF8HwrhjoC10a1fpCiJf07rgatfujcY5zPDrvbBaqTqET0kZZoemCK
SE6Doo/kFjtWJohfFbdJ8j1EMYnOdGcJqB3BRipQbz7XL9NTD/KXgRcZH/6y8Nom4nhv1G4fnUVR
N502Rx8jqz4CsoFrtT99mB3MsY/i8ngGd7JfZO2fQmzcOzz+MgFBDowaXnstHN/OfpUETm3teoAY
XMblVwqt9aS8/VfThT9PRXrvNpkS6gRQblecC0BcPHReW6GdwBG+nruOcfRvPSfrawYPxx7lIRGQ
oyE/fNy+H3zMcHrvhC7aqocOSZ0tkHtGxqp4es8PrAuvKeK+0i3le1ueW+APFWLFOS9zpeJ/5vA8
tXsv89OXTnePelBWXffnhzjnRTGlU6r0j/RmMx45zX5lpfXUVxhdUPmW1xmA9b5x+hsSdK2FhoJ5
h+9O5uXVlIanoLQTJ3/gwXX9qMhiET18bFDg5+mztSh5FB84my46JJsd/YCeWlkEAkqLnndSLXsY
0Lr3jsclNmtjHI5q0+wtph8ilnJV3TF2ogfdZgvYR6jK89y3u8l2Sd4r3Ra0fKUeJ4XSBWQ37Qek
bQH7/KxVBeIg0UJyEZQh/26XKn7A/RRGP2Sm+E+cL46q9wM+LCpjR0TaHsLXrjLqdqQjq+BNHjky
wOALgGrMUGT4OB43YSYwcsTTi52eR1gTsX6DeDdBJvkTDIwGg2yzNCYPvU6vi4jxOS0KN44EGY/v
Pq6efFL5KtTX+jG/S7lnu1q6o3hkCbRIDR5prU4Dh0CF2i8XruPdpMxHwmXJDF4eaa3db2LOcq9S
MqwVe9KsR1UpblDamQ78z0FPPoSlTBDjz4Tr6Ip7r5/Qn6nef35IuP9GQH3hEeX0zqTDKPJBwB/9
Z4+CX5/ZCf8zBlm8Q8UzFPMD0jZgewYIwLgm2UrTBnq7J3JpbJ1Pg4pC6Y/k+74IOxoUSTXzEWN4
ig9YcAxbpkjiBy4bbz07sYRfqIFWf/rv6keYZl35gjyYY/CdT/p4tfeLZK/CueFmzaLxcWlyik6U
CY5GYNird0E2GploHC6hLUM0ZhS0OaVeasj/Nm5cIuapv/w6eS80/m8dbJMJ7aiknrsxhpnJa4aP
k/KMbKelAO9xSJWGh2a7CYu4GfZwVE1dw6QNCMPDZAiC8/77DeWjRAyDskSy5LTiff1NQ8M33sAO
eOTMLz49pNXi27pOuQ69A1o2bdvbZ2JLOV8qgCOFhf4YpV+GLAdTJeNZ98t0yCFBUtPq26Gtk8wz
hpB86Gb5ej8MvNvZwzf07ou/6yQFLjE8QQFqr1Fi9HZe0/gMxNaW65vFaCjTIZXQ4H8YuIbVmBrp
u77s1KvQLwPVgJfUxm1Q3FEuurlINPaRK3GlXDuRDGdtSE/Krvj+d5Y/WTcZEwMEGEGJuj5qfSp5
rWvyUsZvgwZlw3THNb3BMmM0lbqBlMNMmSyS1ip820ZDUGMCHQBsLyBoaHLG4vS4srzeD69UyTHS
Z/U2CidmUFCtS0o6mO2dT4LZF0uypsvdpgYvdBqX1qpqn8V0iGRc52W9deJLpO4D9ivw6Ybj26aM
vZWT6luYTf5U8yLcVJa11Lhx4tF/OZAw7Eciuu2OLbIRST1NW6aEpfVHDv+OBRq33gxx/3mWkRvy
oSh5Vixwe4XF3rpxd1pAMKXDVZ8SRqt8SIffOYF9ciu8EsYjPgFCSfgRQSS4Q3hQLXo9MKLQMuvD
P/CNkz1OGYLsIcxaeLKplLqOVkUsPBP3YNQ16WLO5KesMz4L0IQbJULiGggg59V3HDWDszWMHAeM
zttf6ILqSJIthnRxrql5/IOT9rociLVK3oUrWmWWmlXQSjh5tAPklQF7X9uBo905HtF+nF8+lr8w
3k3NZuEpuOYHM2f3h/nhwrFY0El9Cc91YjVXnx4az0csqofbs7hSHslrnpmRFY3uZSJMSMcxsYZC
DZL5rH//m4Z4049BjMkZpmx9t54hpMXiMiwLo1iJSrkoutWiM2/26vqH53xXaYzVZIiE0mlosYaJ
Fzzz4VKPLNKZdqOH7YqUbuHKImdW68MdSibPieM4vzxvVq90dc+XnZNkKPrCZYHBsLeiOt/NGwEq
ItpgoYpkZZervz44zI/vv7hu0UiKPr6t7zxr1ck9k4d2HR03fUtfy7esnYU4lnV7NMrwRWUWyGfK
II4RjqpQKcKzsAQTGIsxCauesayud26fB78vrHvzCFUs5sQ8686sifw1YI/jQb/7V4dcBZjmTt/a
voRT+vH8U3p8SmecQHbW8TgzXbT+ebpF/kBlp1JQBoT4rW9QoEdNbHSWgSkjZ8/sO9D2tT4qIQoQ
MvZZpkDbO5nKez4S+h4UABFGW475Tnu6bW0EKypSJ6I8XmZBLkiom6qkQD82hwSkqk4ZBNYpfAvM
37I/5wqgZKkq/4Gz0b+RkeFRdAlE30Wis0tvKg9u6Nb6cASltidNkr2JOGM/TrV3fxSUzyoA+Vvy
NH0sWY08sTyE5ty2LuW6uTru5U6WC1cgBWfFXJ0yJ3a0LM6kAL+UwBv5zWeBOL088ts9SKMpr8iC
LmX/nekZsc7/DIb5MCyzOv64ff7U4gdxX/DNZ0y/JhwqTE0PnRoK/ciAj7SX9keUyweC13NQ9o4s
LkmTrzaJ6vTOF+v9FHtkttGZs0xrj+KDsT0FTq4DGSd9VIdlfbsZ9cF+TKiJsYCLYXcnnmE7+SYB
ruUiB3hjjwXqn/up1ZiOZKt1AbBZGUBw7/UDYerWDrGpl5bBDYHBtkDHCuiLNLZIOLqx/hTC63rz
9RZTORjclqw3dwCk9v8PyrFyfSdVwZvf8vXPpGSMGpRppAKMIjZuPhXogpTHkARU9+d/P39ZMVcu
7WEdxEiMpTKOaB5S1ZVCFIXrFENdSRzRwasUALLC1eO8zdTvx9XF6+1K1TvEyj8CH4NWmVcgqp3N
AFfTJPbC6cbnp3z37OMBYdU324w5CtkbwZPhiaO7OmN8QoSDazdpa2zAIEyHst70P2RB0/JLJFts
dtxcaZu9pARXq8MtSsAbOlmpB5rxFCVpGsOXwokkmFRobKbTD/gHY3LPUMoWsDiB3S4ERB7FZyLD
9S/wBMPjpESroPsIiUYPJsBMk4ESR4Eym+Dl+krUUNYQ4MOpZz5eleemmx690KqScFwUAzGvAQuE
XNoM01JieZYwKJi50GuBBfKJgWXkjSh//3FDtF4/dsmdqXMSeAgWn2iYAsQy9pqgguRNwHmYzHW3
sXHD8+lpbLmn78Pf0dUPZ95EcLiiHMNn4LAFJdUCWDYEsIORoSVCWI/SWi5xceYxXCIzCi0EsxEb
eanFJ3yuAZ8gdkQDusB/dKVOuk7kcqIEuZF4MVUNeaIdnt3LgWSzYEx7LhHm/liMzTXcQyFA5BkK
H6L41K3kCdpIfqS64RlR9WwPGdDuNZab3WTK0CoI55Q5xMbIUijnM1PYfqGN6/Mq9AHdIGD+shDv
WsPCcK9POcsaltqaMXMIq7ri0PkbipqdQQv2vQrFE2oyQQUfrXy0JGdQnW+49EwPZtwba27uUz7J
x4QLx67O9eeCziIp+02OIMtLyUsYyapVAQSnfVoMy7+DjXtHtAiHAPf/BQHlTrlcW/vrhZ+YJI6d
EeKmJeChXSoaCm+YBaXbxEo2g7wwplwBdoY/mX1TB+xHx3S5l2r4e4uTCmwZC0+y34rtts8AsZWt
Va8Ror92C/ap2fGSIAmGWXtF5SlgWblhgcZOaA6RHk9OiB6Keh3cOQ1Q1iMnJ86qNjN1rdLIF+5N
nlgwnyGmJYRlC6X9i0JU/qhg3lVKZcd2zpC3igQa3otJOqYQMrF2yn29WF727geA94OzgYr0ZdfT
jPQj7e7d0ovzlVkpxg+rVgPvVJABz1/Ncn60b98JZ5YVvd0suEMWPF/kVHnsVf95D4IophdSkp3x
32WJ6F+EOIX0aYT/qsVmPoLI8Up316+dPkDjCE3BaoYt5mXNgEM8dm96Z5Dte+jPxw47Gv5ZvTdA
Dbwp64cJExds0bDjPbYNsp5gdSc/TPC9xEOR+O3RCxSoKQSPL+w3FoF5t34/VYukjyKYfExG95Hw
ZNau+y0I6JF8IP4ox5zkl2kwYdCu0JnG7XImx6NIfRn4VnoFvO9f8QfMRBGVJXYDlWTeGZL5REiF
kG8S8D9ViMiW1HWOL7mzgvbUVKYfD4K1idiqObSzjnqxLWTk0FFa3Q9ZXxoRrNVrjRzblqgKhoZV
+1lgkH/AUyq66mDMTRD/XERTT5n4FqKhKbG6+IuyT67xXQTpUVaJ5qEKkIBLPNuHnjoZgwjfWQ77
nNa2iDYp/QWdxA5CTGIf+n2ai5C7X0zmIFrmKfDs4nTQgkjCCaswUdOZSSVWuaZlFkFxvFxdKsw1
T3uJJhKDtJ3PVeiC7lzX4z0Jj9vRPysmAeZ6nLJFS7FYFD7ZfyvfINnJxffdZrBy1+xOb9Zog0EQ
5PwhZRZBnazcCB/4bBn97TCIs+K5dnWjr0Nag3kIJzL0I3lBoE3ySUZx2cnfE446KRO5MQXKPRRu
rbMq/5F6qrfeCLqwNNDgCKU+hmJhWa5TmaYcXnO8zUMVJl5ZqmtkH3kz3IkHMDINjKEJTSI3P9DH
FIdMVkbZ7zysRBKxI/ycq1cOKVj9uV/c8R3BRYNNdoIvdoviwqiNbSfIHmTqt0NhPLNMmSlivdfJ
1i1di265T/qTH51b1glfbl6o2aKabhs2gRUjIPfPHwzTfn0AYlc3YufZtFyHdj4NRaMfC1qLfh4m
vT3MEPV1j7ex9DEWmE0Y/hUYuhBBD72IZf6gBKsCQCl7gELk17MJXBLNKkrfl0MG/H8NKyGiWPR6
xg6sajojoguT9Lz4EdzDP48PFsVIEhR0PWwSgjue0HwhzGkgy9q6+CHMOP0a9o4aYVwAOTMACSuu
7ig70mjfp5T0qrkwYmJwU3XcYkPZmD7mhQIVdcJbkq7khoYH2XM788iC20ujkzPbWYr1cN0rdPmg
8qoQ3cG4SMIGeIMIvnwuuwKoShlYPgS8eiZJOmIJV225pxDoQoKRJo7nQG3GznjfREoetVIc/0WV
wBwGN6Bmvy4NG88mJfCN177v3a97ZbJ2D3DyTvA2s8mmAoPfd7Xj0aJLjoB9nMy+Yt2RcYIKIcFR
9040X8cpMLat1zvdMTpmKf0YlQFb2F0vgDn8L6KOj/nCLmIXUiIabRJc9Oj53acQoEeP72i9H3kF
43UG5YIlit2uU/9Wc3Ra95LOMQVz7WcWO2ik4s+hQhrAsXtGW7TUrOVjjKnhGFEahdk46nPq+5jG
cG7Zoe21Hu/YySa1ZdS8sv6OAXMoazVcWfr5BKDD7kZXnYu76T2v1qQ8HT6h56dusmq5/NJbcHqD
6Kl/xOkpG/STPRTnb5U7JRXpNZS9yJj5XlGjd8L8ptWZmP8oxf5+Kb/j6nVbr1IjAZfygLcb+ZvX
bcBAbotmgKR9mCn/WhQRPhEAUCs7VIm2+Ag8QNj6ixNQG/1IddT4Nv+hCNaTNRKjZffBduko84oM
wDc9VYNTlXfEabzZahB9CPLX+U9zN/S7x2o+9Hafou1q54dB/WOisrVB0Lv6WSEYN4DuJQIKC729
Lyu8uCq2D2CBTwlsVF7ljGRGKzPxicEEhLEu4Gcl9JEeQqDJuXk+EXGDQ9T5L5lN2WsuJFwWxBKF
yKD5LkSl3CupW2XUbvmRaPKbhlJ4LVyyk9v5+3e/W8Vc+6Sk7ETZrnfFQq1pWmoIvnBQVl5cIk8r
KoPIDeNVYhbzmo8KH2VQMB6BsS/meGu9BWqfSRbxOls8vj9XCFzYDoJ36saMoFgRHS3jMUtyDS2+
WlgUYjqkoDk6oGBublXBla/xNSkwxbSewFhJZgbnsVDUt/9wxS/g02GWDa4V9cb0HRthz7rYlDCy
T1eWTMamWGPq0XbbgRM8nM3SF7ogcWhxOF+UxwYVrV+dBcnC9X5qkm3HjUlKzRAnsx1/JP01AcaC
L/PwFt070PVk/Fee2I4RhrC0AnJk3FQUrXe8+RN/b8gtkiedFMOmYZ+OFw2KrZ9jzpClGPjN8t44
zlDDSqlOe/QTfmR7fxjFvE7M0PkU+rpdqCzpn4vWjO2Luy8WuWbfLr705CrslUt/5QjvgRXJqQYM
BoVN+FBryNmUDvty301eccQ+T0v5qbBys1Hq+sMpCVFx3/OevAQjN2MJdX+KpUCCJgcPfj+PhdOd
lZhPbDquIJ2eiRD7aQcVNHh7xa5LpM1VszmBM7FhKNZa35zkXDFJUk2M9dFqhYFcwTK+gSUMEPMb
TgK+MlX9ooVQHKBefvdM7KFB9LtUzOo4vBT7ZNjWPjmF9aP7rJFoG8JYBpBjpNeil8HvkGbNA0Cb
W7sN6fTjJBv/MuQtNs3zuKHa+pNh6oKKIJ5XelvEJinoEjJ5nDF1GmYrxLWCVsBCLUpLC2N0e/4r
0gJlAXP8p4oVFaG/9KTe54uG2lkCLjO4XA0VcXMlqr+GozE259QU8IS5rSNwr/5tKTfaql2kqPdf
DRi5CIvC6x2TKpgC2aykKppGyolUc1xIPpWK7xdAjEnNA24Fy/9MQWp1iIo/nf1Z2XnwZnN2+nU0
H+9imPZPoNfrq41CsUGY7QvuwOuJRk31cW/rbr8zKrKcPGnnMoWbGZelHZ3tiMPtKMBPVbxTOwvy
My7iL7WswKt0xKeEceUbevK0q9yK98u2WIQi3mEvIxrnTLsuYG0xbSlFRszhTZcKqB4ysto6JaI9
bYP2Ga27TqEQh0DI7T0Gl7ETwXDuj1JEwt5M7Md597HW8VR47cp70Wjb36ZCZPRG1rGjf9GTC+9Z
YPWjTAPQClEq9w+TsDBE59+Jb0jbbJMmGhLr6kv5wQYiMr8LrUwh6kyu+APIDF19kxWgvEaWHgxT
+VesVDfrsqSTON0ENOaP7rjDlRaa40iu2/KcTbv8qGKs3nF5yIAVPcbCd17SAXnQ9P5n/ysgXYtk
qlJn1+cdEeZ4FXxp9WZFeYmxzOnk63SaM/vhwTY+wd35NeNHwDQZAZWKD0DB0QCkj918Xj2sRHlS
pQVmfJAZSC8v3iLwGSbYm39L/D0BkJl6EfG1iyCDx0rs7c0hm4a9mjKq8LSNVn91n5rlV0nHt7vY
vDA1YD2jvQCunmLQXy92QtLUg6v5BUOZUo6ADctIkFCNHBgATeHbW4/1lVaNkw5Wmd0IVJc4ihO9
CRJlCxsGNy+MZX2R7GZwBg+iGvz27tTkWmhXN2P8sM9/otM528k2iLGW7+mlbArtwrXtiMix7AJ9
1uT/zdBsXyJ8NqU4qsvt3pLFBo8Mnea7LOdohxZ88eDCA3GI9vIu7vtEg2DRz8pqaUZQG7/cXl6f
ZpHyWOnLnxlCymUDf0SbFO6LwE6RduSF+FTULXdIs2A69D+wqA+xaHkjKb29K6Qcb75TNBEpYx8Z
7PYr+R2kak/bpa21ZyWGSvGzy9e5WfZy7/hjbI/WTJjrL/7W+CXfbw8HzC9n8tEgqSAXdaj+ZKmr
5AlD2PBEqvlkaPEd9vKfoFNMcXL3X9DF0gVjTTTDB/TqxcPmVhCIFdRYCVCZQc/dUSwFy6Av37V4
2i0whrBYZz7UBlAx4pewXhk9hSf/CGMFe+l/k//0aXyP6k6NR8uTwrHDCc6yRYUKDoXogGQ6eHtK
82b6ES9oJ7llCYYUFaPvWKZfO+n31+9YYMqJ2X9qJOdhp/JhqnZrom/oftQFCv2h6Qc5Ltnsccg7
kaZrbLAA8XyPG7OYBN6pVddUB7y+3EdkU0O2XaIBUlzrult5TtcPPnPtWqwrCHLa8Lx4U1Lde2In
rZGenXSR51cZOY8UYagI1R3pDkc50BgbqjmYJTd0YpYDpjSHnscSOCc6BLtdVF/mi8uc5AkqcOuG
lRSXAt6kH5IPvdKDiAihydeqBy5+kfbm3GnUcmbBO5inwX+5h118RabYKmffbazUzA6eVKL8trOk
enYKzxUmuLKz57QMLSaewijZ2H9QnJI2YrncygxHD+qcZSVAThpsaNhODlx7d7Mvd73VaML4/F5G
uc//EP33bVNRdEmYi2dyJDHNY8Q+B6Kkmv743fwE9HiBSZz2xY0FQAtM6rgGY0bWT0TB3Ail+SXd
MBJo6aTZyG02pmgpXMjbe54DNPvkeW5paFOi6VSrDmVT6oRzjCWpMZmHl3siybCccGJ1yrtf9qKN
kr4dsFyhwhJ7W9GLRsnJacscZ549Kr4YrufRQDxNHmaevp+q9A/HHc0QZCNZglrim6xosUHgaVrj
HeVB6Rx76sTs3yEMz2a/pbXc0WfKesDkn2Ie9Wo08HkFbwwrRmBKpRfGX44Hl8WdPATy9qY1Uy28
sLAw0YtFI8W/puS3vgduLw/SE5/8grvVy9oc0KzwJzqt/SfTIuh3HPakQ017RharsH/XbD+KYq1Y
xzui+fZLHFkMtcOGjM1nGnuvFtqC7JNiXzsNVCfnilDTvYeyexr6aDaFmOXKKiMTp/fBSAohj58U
6AYTKQOpc9e9poVSbwijGH4mH2yXKtVi3x41InRw9v+F86+HtFi2Pj4tf/XJEW4Yaft21TKC1mzr
ykHCIy8jHoNOOnscrNn+DG71ATSVhI+CHoMJXZN1ghCDZGkCO8qQMfechUXYPXnq9qIcprIKYm74
Bte4c2MkJ/cOjibonTxUfeOvUff/18sCyYBxRANnDAsIyAIUTjZGN0WORWeQhx4Dm6/T8QFbbQqL
aQiiodKoxXlVrlyrhi8CPUvGmYcc0WW73j0f3Sbobe3OruCK6lvMaOh3nV7+QcXr+iM39hF/F6NR
2QyulRlgE+TLr2asJc7W5hkq2jornm3MBsdvlaRb7ypWmWWUkDrOaoGAJWik5O0kYALBjiHj62JL
+UjZ1+tYgCwkcgYX4Nss6Z4o85QghheCPr0xTIw0RQAt2f8FKLkylB+7wUlJx4q4cpMnjuI/ZvIu
G67bvCw6ZlRKVVuVXLNDB1GCNqohId3HXkWQ9V5oi5Iy686Ik/sHEmqGP+HJVhJJ3lcvisfu+Sz0
TZx0QEQVg0llfHsC9qqKD6amx7HQgsl4HXCubv22Lgv1EboEN9KvUdaH4eQ04lHU8IbibI7QzDj2
eaXw6QIAusxO8xQBFnWUYvCi8Yj1M52MiGG1EHgWhuZvnWg3NLSF2d32Lbn1ekyEgK0beJJ2rRRt
cmiXRNXagrX4bQzDErq/NP6EcPr318PsHKBVjlHxOxlTVLOf5KW7n6MLYKpoZeLha7kcgEV4ERbf
64viXYA+X1GR5lUnWobXyFIRSijTMia+RB991I65ckR0UJvUkOwRZcmVyZBelAomk4LJxzIM+ffh
23RqEHIBRsYWFAIIrHRf6luCtu0Xm9bdxNMtG2vKr+K+lJ4W+rDRLsxtinv6CknQ69FnwgJR+3hm
gyAtMtWRFA13hlo1jUwj68dzDXrGYZJcuZc0zbjkZQChTN3DZNSR2YaN1q7Rsd66S8tmxLRRmLVn
4jgRsvHUxVpWj2Esh6ceQXdWeP7HD5FQHUZtnAf0BlbHjBXNsGEHYOMVf3rMuj0SkTyYhyp40Pzc
tIi5a4TeRtS0djUIZOt2XxQLEgTyhUSaJQn1BjQzolDnY4+h1zqHXrCbdI8H17ZoT0uiVZ7QzmJD
/xRHQp4bv6dGnMkERzO2fhh+SR5Buhr7JYXiPEGrx1Qf1fWaJwQ8AWvhzb+t2J1PZFNn4bpwP8Pl
p/KZjAZ7wKdpeDiHM46a/XiEIfdT8R4UbgnTYzegb+VsHwQXHqtuIWtZfo58kQKGy4COCypqPKlg
upbhPWR4INbet5odqqaFoJzeAzDkWtLJOTNcz63ur5bR5wB+FUaSpq4fdU5dMjyN8ya6rtjDGbqY
YZ8cHzDJDHOhblm4OVUO5FmReGxOxLwRqNC/RpXrPHhWHwlBZ/S4xkfvn+SfIzpz4wyaNBXoEzXS
joIqdRoPSEeIAY1aqMTbUeLYEQswCF/Jmalc6H1wNIYaEqLHag0JbSfU2RDh+xYDm9Twyj+Rvret
cUk2w8j550FCw+qeVnF7HbAeo6EaV0S0mtm4F1atcsJgDEzZwknIg+gvQDBWOU8NmcSimmBa/m/9
ZZxb1KUZTyUZqm1lHCQ3sDwF5KtmVBhojxGvGH4qI7oyI6J+VhHut4ZKdY6y+fdu1MR+um0lxtLf
zJ3jQPHXgYiBHd60cIqfSG2KLkHdFeUHszDKHV/MiZXg4jhjBFu3AWU0zTsxAU/+pnqMsTQybLzd
yQUY3Tfn4u9M/smOvPcbnh+RG7GRiwvmAfIkAPTalw+6xbvF5ZFAhsBcaeFFVLsMFpisqI/Fy0pz
MFallfvTTyQJqpGxXinBFmHP70ci0WSQKTfnfYGFDQJFED5AMv15mV+3B1kk+NgpMhRC+kpo7kmy
zB6zyxDfZAZXnMibt7nmqwtz4w6SZyDAakDcNypcswpsfi++BmLdjt0rLKBZbfoC49eRZI10U+oR
xG0c9aHJwTwP20mxHOiK/V0vBbkgnYRZW8IwLwQvHU/i0JvJWOmvyicN023u+twv6UHQPVgUuBi9
c3w1+RRcty3XjsFFdT5OHnqkfMkHf36BzpU4z6wSjefNHZ1RCFdpBFK+kLabOm9VgxIW5jdUUxlu
Wk4Ef8pj+b4u4AE9fAWVfXtSo12SPHXb5Le3BtDORGQf9udDrDAadyTIdSNFt1DhVSJlc2Csm8XM
CUlOj4CoMqxv3CUXVaMctev6CExzKG6Hl1kdwIVDscLbIge5EQd+NhYiQH1Lh/huDizMVm0GPCn3
VOs/QOHG/wMwruUT4k2GTtpshuHJojAH3AxaTEppbnc90thdTCTIvsR50Y4aeNhHKpqeKuiRq4z/
s0kV6eUU0cDnwzU8A+B7/AIB826Zy8im+Jd81pnLthhroreIvvbFvNorun4rZSw6qoGAhnfl+BAl
IK4vr4/hwYoLLtxyUPs2MqKmbLynDihMuDvruQVu6zbWRXWZ9atV67CQm+Ai8H+tiqTYKmiaBD7v
vtklKqq7CDV1pfaLUpvKHp7R8qTKCyjP0hdpZBTHb8t0w+BJk0ODdWNuw6trhjlunpUTJmU9z1wn
3RCQuUbig1ikFPiVk3STTtExpqopjma40sOEC8Pq50VzZLtpggBs6MKjRewA40yzoDthAqeelUC1
94u0FQ/nqN2ZSvLOLMepsInsYAwUbZy4ihZYFTizf4AKSdgwfho2QWExqmKKelIPgmyQISrUkocG
09D9ue02lUoxEngX1yOMFo127qCkZv/y4ez6XPwHVu2uXV4IeDJW5a57Hp1maLN6WXez6Z0mYsed
yveJQUoTex0sv1LGdR4Y4Tfsvdw+Bxga3AlOOiGFBDvq0JvSR/72Dx37T8xv3UYabYBXJ9BeG3p2
+t27aE5cQCIyBXHqtvl53XWhHWdcremDgrMDMRQipHMVsl38OB/tYmAAX42sNm7U/WRgeWy/8fXt
LgZrCjSxwGwdtVpShxv8Ir3btiG/2aoTKmn6zDL+cZ3edPDyJe4sufiaHeP1ISW2gvZifUVtpgO8
Um75CDEgWAsHTNHJtLBRd4TFQPd3aV18QVP21febzEIH6hLF9aACZSC0gkxjpnJvb/kUd1y1V2LE
PtKfEa+xUw2TI1VuBCnYYwv1otfPOBw23i3JfbvyNbjzsoV+B1+G6KD9wMEBxQwuf37uSQzD8ClN
rBjDFpZfZj9ntK1NeLMJvigmF/dt1NvCS4Hzw7fXxQ5GKTDJPXzSemjSmhDE0sA1zgcoaBjy1jKB
eSMZjW1jcc7SUg16e3gKv0zg0BgESGh1WGPAuaLoML4KvFF2t1WbHa6mmmgmiC019C/gV2NdIbe9
eKNn305N34h2veqiNvihwLb4CPyd769pNkr/ALng6U/RNnO1ye71ej+lv71odGeC9q5h8oOLAn2n
MBduuJoCTifMOB5HO23gr6tOTWjCpXHNnPSHIyA2/ckLC4S91pL7tPzQSeFcrxGUlgq11HZ3gWow
QRu1WMaec8NQE48aM0K27cIbPOh3kjF5RLNudjGtA9NBm2VRLYsJHyWQ6njzV+JR47PK4p6mwI7H
w1DHsftFEcNJ/htQhbVtEpIlsENBg+4ym7PyyOQwdwmyKGreHGtc6T5xzxLDzquW293CWKXkIdnM
oZIyIZwcbFWDwQTKQAqlxYtUP+bicwnNOpDtxd0BKZgP/HZhqcVXRnoGiDflePV/czPOKfNjIQR1
UMwTJIKa1uVQKUCgHsWxCoqkTItObvXARyZtejM5PRGvw3TRJgvq3voNf5MxctFXZQ5en+quOPhU
76GYVv88cvdjfJXqcFsfoYtZO0GWcrBBDjvie8z538xkIoSTTcojgzBt15jVoJKqt/FoXHGhTiVW
ikjBkcatbenJkd6dFvEV4psBblHc3JlO7hRypt0Zc+rHE23ZehwqEGpPxFQtNjEgkX1LZDe9+E9E
Dfct64bKFRQN0h7OsRNmOy1P4P7DFDvdntueZvjrihIsYi714jPH547MR1dh4iDUi2htN7GW20Sw
QWR9PNa0UsXqR8FiRdm53sPO/+03+Gt9b2PZ/QunFYsS/LJvRbnosc8ipYejGWcscLHrJApJXTKo
OTr65M+vHp589UDu6IkEtjGHrh4TGx3kyzcPZF8Yx3dOXwJgqs/vMLG5kIsX7Sq1o9Ps0/p9x89v
YSFr7L9IIsNXT+3dvNprqiqVp0IZUuVcFcj4o8cD7vACtNVO4CsfNfmBZUwP0+I/whB5Fi7UHYfx
rZX15j8hH2nGtNuDyPqkussczHmMdh4mr1DGihgKcwAY13PUK4Qpyj6HykES/yZcjFJlWh/+p3h4
7zcp+SjbiUeVxu8uic7JO9UcE7NSgosY8JWvqQlhSSM6CglQkG3WmQ0mCHUg+hx7bmsO03eRUUd5
BkR6yB6BmRgsvmR2Nz2MH1L2bFxPtrlX3e6++LN9lewQlFlt/ZRi3nSp00azjmoklQvfACT1pPPa
BE99xP5R5ntv1xbXRDmxvJ89QzwBus5BSdImobUKRq/zr13ltpwiSmb6py3yNVT11FaVAUGgyaXh
pV+pgAnTMyk1gP/RmCNTeQbAE0hxd9Tv7brvzBerOTtkofoFig74lGb3yv5JB//mI9l+sOPfUVQT
EXJGmCAn7qC5j63DWgPiqHNFEh0aqYAhQx5sFZgy7oVqZ1B5XNX/3ufsayjJKJ+PMXeZsQRSoJZG
40YeErFowmr3mET1FtvVfR8Tinv9BaGHmMlX30eVIXhhOf8SJHO9BGLL2SHlwd0vbyAjUg20thKN
e5uaaeHyRIFIPCCChPOoolSAlJuu4ShTf5MOCt4WS+CdSAIrgjUSCvvafLAehIUiBgAV5Q1Klexv
YCEGH/MiOFBCyz5zPFRLvUnxMSWhcYTWqB58TiaiudkJqFx9tH3xgRI4ZtWt4tF4FB7gB9TtcQs8
6l/mcRJ9DYsqaoNaE5S6VaRfBp39+0P5n3YLoXSI/X0UdG/YgCZGB0Ebhrzwv3FI5oWipblXeD5E
eE2Ms+M/k6kOCnxlipFug4BblEs/kEzKuLmqfo5cZt+Su6qaHLGg1ehhKKAHFkKxUSASxOdV0v8Q
2Jjt4KiSSLTKH5f3w8MMJ/pm6CSf2IuMmVt+4mW+Y6regb2RvUITW0kP6wkHSDZpBNszvN2s+5FK
U2rwGWKG4LdQvbaH7q3DooUjkqdWR7sFmBo4ai1XvJh1QYk5WgPIypDT/tuMpqsaesUkdqju+mYa
eTf2IInygbbmULs+zkzn9kBxAsHb4GLBzleiz63uSdkBsh7vX9HCCdqPx7x7vglIWyAIH7dIbi6u
NbFChUaX7WK9858Jy8g8fI7BlNK29JgjJ95syhteQZWiEvmCVXrlf9vr0gGGspAEGwpTERRHq7Wq
Xi8LCMs+UpVGI07SNFaq/cykyEYzEcwLzHe7JsfwznAwEf09iNXFonxUytyLNYQF4sCy9qVMjul6
lNXlO/Sp+W5cXiojZaFTkHAuCqZ1gW+936HlXA3C5C7sE+v0QInszRVAHQ2PFM+ErQSA522mJ8hm
baYY3RL4iEQe7BWwBk8WApfgO00A87rE4/BTh/80D4Xt5By/T4WHuVQA1VZigyPRVSOejFmCaKj6
JFbXICh71W5CqND7Xz3UazOog+lqpwfx7PKBUvAmdqQ8r3VFwZJUtjRdruDOLw1mZqZM0ncfe7S3
a7Z2GvLyFHqL/J70RkTZarWHDgqBkPwkI92TnSmRLiQFHkDEGVJH2B9+XogYyF56ukI4N+uwAnU3
3dgUPXj8Mg74jOZdWB5TMd9c4ZtTDTCkCwWXXU+pMQgRvcE7/d6ZGqNu1DmzkpJayAoDC/9zxMOt
4RS0mSxr+7LM6MOPpZ8bEZFiB7uRhTcc8yJ1zdMaGO/pysyoTb0qUaqe8HNYAIh0jv0eCpyR4JTa
B/lJxKbvrcLGA3xuf4qKyndDs0xO9Rdhpkz6m5k5W63Hm1Knu/4GI6fA0lR+ewS/54fJ7LkL+zU5
FLi8ah2wdcRQj0ZeBHjaGVChNYJCKECATpNkaJDX2i1bCIhW4lvIgXZzQOcM/QPtnV9u7fnJVk5b
id3pxOQGf3lhWTvd+rQEPPK9dW8c7q8+inFQBt5xG61WzTTY5ha6cs0gzBnK79mPnpzypcCXJVLg
WtBCOL0VqLZ3jz4kGQSUfTgMcfFc5NJ3QOzUTH9gNgbP+ohDZ/WA/w4rQfChMkol4ZMWc4nt/6gy
y1Y7X2UERpY95kflBTT5Qay35g6JFyh9KgAZXgU2nHDdVjbJBLUIoX78Ko+gSgg733lm61TYQVKL
Ef5tKM1ILafsm4GQ+eJNbre/0AOYUPwx8lYpabbSfJ8IANl/6TtHlaN1IEbZgk4D+oHYrSEnlGae
ftIuWOej/Xv93je65owWnoUwv8na1B/VsGYUlyENwAt4mFqD+X+wCTnpPRRjYKF1WDP8RoIdPUE5
3r6uuDqAW1cVdaQ8316jFFF43TuG6A/L0i601E6S0oozz6r3tQPvzoj5lp4zgt7inQOTk7Vv1uzW
uDrboUIdhxDRDTfCaspi3A+K2fCiRWRbxGe34GIz6T4JmA+ojjOCEG9Ijc6Eltr6jE4iSWsnxQ6J
KPxLTzrOquYRMPPK2Y9inF/NAWRLRGmB+pzvj4Il4hfWcLvg32EEGIf/10wIGnxtA3JGwtm8ofNS
YjVBGljvKsC0H3EA1wQkBinJaic55i+C/pUXfTu9/JwRffeG0z0VmVQs4940su+ff4Khc0bVLlkk
OtVKE1KWQi0ruOMF8WfVJb+vFJoZQmw9RNKsLtTsUX7cu+/ZOF1I3bcOy6tC14uq2qRawoXN76JM
30YXncFHzr9hN5K7+cQkE1JYO+efgdV/UMcaDh4LNaam5NV7SMGLko22PXqbC41RkMek0Q2t+nGs
WX5okhDYBXnpe3aqnEol8m1Lxo5+olUGJcX/FJ9/Ure3Tvqi4QueMMyxLq/fxGbHRwCg06SJUavu
X14KpKqtA9StEWHxc5+P7DNz7RhXnkF1pmMuChtzpbMVsPwzZIoD8KMGB2FAncUg8VnEaplWQ4xw
blNqXus/pv+6/OXzHMXaltHaCnI9sLpbRMinYkpfeb4tgAByeb6xnWw2OSoXjTvGWXuDPbZw2QRt
iV8QWP5Kj36bqirZZlNnceRaU2Dqxp+effEeVqM8f2xk20f8m3jezwj9jjy/RsqvcZ++OSP8dcw4
waUaR9T67qAj9hvsbNT40b/+f9rwq3vTshIdP8QsXFj4gtyoqJzUe+AN+hGl2w4vEaEH5db78oJ3
IBYfPlSP+2ID6r/dQy73s4Z9HKEdUsW0F02rHPEBj3uyU2pXomtYJls1rEubCqWVoJQNmO2iceUG
FpP5FDYjRRhfod6CbRBu3OzH+SgGhcXKD7LkwktqSlUefMmFea2xXBT+d6+hjuP/WCvQBb4f4uuT
rW0IjDmgyGGHjOop+5fIXRJt7kHrrmR0HmD0KQql9EypiBtPGJJboTCNKfs5NRBsygbBkCFOJkDx
WwpLaoqEOu0e2LY5g5NlpxJUOfWyJ7LtUqIKOD/DHcofgMopckiRS6tLE9bd5KumNL3T8h+ftx4G
3lJlRWlvPMMonHkVjcdw1/K1Xt7fJ3USX7IiCDOeJeKXVMZXPH8iebdOhmgzjVtBkSLXpfMv3SE+
EbWpp7Wi5D4hW00kFbtqeIcRp3KZhaQ20HZ8VpncxzvHi71vJSvR7YN4v5CbbmINK7Pc5mEbYhio
ZMCbwG0A7iAIlDQwAocdNVHUFoSJyfISbi5eIQ9WwD4McC/aLfxurU5C852Mw8XBrkN3C3z+Up7W
DtPw278OnwjVqySW7+/MNqqiOHsr0Q0kWRl+YtaQp+2PjSA8HBo6W+WetsZT/ZOqwhrAVfwcd2gC
w7FTgDvysGatJdPUSEIJYDvZ51GNpq9/TT5JuGGaiT4xY7IykGVgPgPHLtLrZTIgYbWygrKyI7E2
pccJjMpLx/XkPP8lguC7+vJ5vAR55n5WsEaHmzkwsGgV2g0ISqLEp4V2YP5t9uO/9F1qAaPLATKk
+8bmHNC+IQXPE3IyKpzjIXAaLf77r9+O3v4GbLpcRMhNJJQH70vwKR7wtFdCzawCaBkhe6BhIJoO
wAYiKDutZuV2ZmkiUKOMZopV9Z1xeg3bn+UDHQ0W0O73NcuE7N2/RP9Xtwv6k3xJGEHwKpYp7TwE
/4JPubuiqJ65Oaen0DgACmxPZosoovn9RY/cKThLy5KQifziX11ULGZlhlnclOllik/0YWyeYb40
h4vRPs7QQc6W97ph/V4cErxjE7o+kgXZ9NOGJCepCNytbzkhlXetyuFFssYKciiems/gH93/L5uR
ejG24tut/uSs+SKmMP0LDd6N+eUm/puwIuXleyH2WJvchZ5BuebI/0Kb3K5HyljL2S1bXe6j1rtG
UJ/jvG0wbgj3s4PWDRuIVBBsoGHb3TXdBg0bzCsqP6J8dRU45tKzHYrDQ6OWsn9R3iEaVJ8HOTFh
TzlzjKDJVz7a+7cUUSzqxYELIi3Yjm3cx4NioTg/uCsS4HWvXcI+8bBhO+svTqvr5ABQ2GM9wPKd
/04XPYeTFfb/0vRkIeS8xRsbXaZPvE6myYBigPEw/uVbs5G/ZOV+D4LRFHhAilYCHNALpXm/3lQA
3lmItDRES1pzsEcUBIm3Phe5ptLN0NLQ2M1TM6MFAtPUKyBkic7EzdfAtkdnd2OwF/6B1sBsBQaV
WDpNdi8k6VJEU3l8KSrRffoIYNrCODPuHUH0H9kTxehQ6tI1gKduo435qlfuchqlz9P1NoFtXZeh
gutM5nyDibbjdhCUw/b4UqOdAiG/MN29bC4kPYaAXrmDDo3baGPyjGTGT2K1PqPbA9xpzA5nJj6s
cZ9caaEAi51TJZz8gS62nP++GsKIU0/0d3mawnTXeKNX2N+FIEkKNY7RwYgZEznHW82ML4XT0IJ+
cNhVlopp1xv3otcjXi6z2Rqryf21PGtOGFQGO/sfY25Ag5X/dBwWBSsyQ9FvYUzF8i0pmT+aDXOC
J4rKZcZEWjpDWkvyQFSsOIzu4yMXTwx+9L5mNBSLhIGIsNlaPzGX8piZRrl1d60AclARpp1MKpvX
uEIZPAtQn83Y4f7PFJd0kP2mqSL2XFAlOo9jd+S8P2OXdWl6m0xDCzC3ezA2SIcgRmcfti5pjH3B
UsVwu+OVKOw0XwcXxG0tDMYdlf+DAIo6YKftKWWml5N3ZHT1bcXLt37zqnyNec1v8m27R7nz/Xf+
rk2qRDRW+CockrMrtJo6H0mTryT5saGRzX3DERwVTOSbTFUFivIOpyYptDQ+Jeil8LJNbhw9m1Xe
xvsF7TyefOYWKmKcE56Q1PhaBt/KZOheiSfMUiy1bQTCoUDxYj0+f+TnI86ebz7wkGKuzlcrWRnF
/IsixcI75iE4V/NYComewH0Dn5wRG4KHOggm2xNMNFizU9ls65TpjAZvNxGXltoKz+z0Yz74yue5
Nb58KenayaY6HCSTVm1+faWGCs+wWhUCm1XxN318PTfLBwevu7Hg/U6gDeLiZAV8IAmLs43/qkkB
Ge/rpP3kpA9X3aEWrA5CAT3U+rGezqyQCnJxXzHKetbgZjT+3BklmGS+Wtha5poRXn1q1SQyygTp
/Si62b1uaGTw/kFNGCbgWlmdZrW/o0L4JcXs99/gO6O/xyIPKckOFloR7LbtWcskLWpkXu3xujZ9
aOHVhbafsqG3xzOxDg3SqzcXznJvgfZo15tmqTt04en3Fq97gbxPccifsNfO9IXKLUAt3CWdWAqp
BCufKZnkpqiA5X/maaUlxE+qa8eS4zlW3ZgNIKd1czZTjx6oRjjJ0IVs4YWVz3bhLM7Oyu3+fVVS
YquyeeNthdeGn8H9i1+FguBa6TEQL4PNjKuNSvdx1vFzUZ5rkA4K1T/I4DnlHsHqOzZ1RcoYlbJE
2ba8Pb6qTc9Mw+CQjMOQ9rc6TMR44gNNwuBD7wA2/D2zHcQwdkyFyK/rAiPbrC7qOun7tVN2DG/D
y3bNaa1ftKnmTQCL3UqkMaIdPmNf1qk8CVQH801TIC0qI39h9Vf+0EYA95YG1In92oIvvOBjg1t2
iVM200xTfRpG26sk9gHwpcLZC5zeCPl3bweM0jprPpA9/TO72R8/+9H+wmuC83lwHuIXvy+jIDVU
7lZJ8eY5gBapOK8aV4Jbyt3SOXDcAwU7cO/y9Ehk8q8TRq0uyfCvlpdy0mqsmUOdYorOcxdsYma9
McHBz/Tz6BvWLz/M2Woj05BomJ66YnlDi6w7j6cPlCDmAWvxRzjfuc7REJcxZKdf/fq6N9xJ/jiv
zf7PZT7Khh3o1VRseQW6bFxLbDGDIg1em8ZlUegt5vDD2XX+3MzTa6NCZj0BKVGL9N1/oAfY/65C
8cnZuz8bKRKOOF+kCTjc81pBalWBy7eEPvb6T2OHYpJfwhvukwFsVA5GckMnTMcb5tx9Bny/O5KO
4pL6sHY8VUlH3Wj4AgL30CbRpJ7wcqwOz6AB+i4n63WMXzKEdRQj8W5YfLgILvQteI8P2+7aSS4Z
+22t2HvB43l02RGzVFI/0mU7nvx/JCZb7wevqbZcRKACqpaWvdTCqQWKc3O7gz0niedHzyq3jnTd
nQfeW3p6Ss2KNw5ULsA06e9Ksijnjb2Xid/uMgTDKc8aCRH9RyQkdHh/3Ze6qoWA0wcbd/5I72D4
7VBLWulvxOSf9xRaJk4n8WZ3Lix68coKgGgFK+REYnBwl6ROexIZwL/nOVs2F9iOtfN3xzQZJE/B
6p7Mk/ftqmohdm1w2kI6apV965UvuBoQMOKEfTRE72L7Dedail7qSjGiZlkiNirpxKSvOfMp1Uj2
ty/xe9AWg854YndEu9V9n/u2v5eyHP3NkOJSkPfW+3oTzop6uzqu+N7gPuQE+epeWz3DwgvphDpu
ZI7zcBD7csz2c/8yv+TwtiiFXzAo6lhCoWJ0v/EAVWR63S9qPT7Fu3pwiE/oLvMd5ChRnPwvLDL8
bwHdYkFJEzDq+dGpiUug/PUNGqj9wN/lfAaFMts8e+esi+WetSQszxlIHf07B0EhPVPmLiUWYmA1
baYoe6eGxZfys92ZvGGNK4ihb0qyJ3IESoKu8P1mlw7mxClxiql9kOTp1YJHDmuBFAyxKZiVTo5d
FCS+YeQ4PYodKbhVOeHFKuAxdajHVnS9tnKP039O5h9DXBaDeILELRlcdMx5S/V84Rc3NaNq52qj
ZQ60Q90IMfHO3ECQGRHq4GliqnEg3+3flQiM/mslpq7z2LvTHju17dplZYbL25QqW13+jNgCa5Kn
cRL9Cm7NkE4vvKRY+hIhkvALV3PsPEHzgLxooUb6ufq1tIiWTPswlFy6UmkiFB01U1gbtaNBcSGV
KKDhFV5uFoPIHBiEMUjz8iEb2Fuv175u6q0FQ6aKaHB8+Y6nqKVXkg8KcWzv/vZR8WhLJRQSMxuz
5s/JoOK8RKFJ6BmxtzmUNPqHBgueHA3J0Jpxa8W2eCyrTs0JlTRsnyvvCN6qeKs4EYLmCBmdv7pL
PFikEFkjn9pAp5XqyXOfHiQe5kMTMTf4b+0XVLdS53jTrqLGgm7oPSjKhxPBTFxTKkyC9FiughRN
4H3M16fxYskePACC0P8DNtG459kQ0OM+UsFBXKc5Bw9t9iPmJ1hyJwIh0qNfaqxaIaJKSIKpt2AM
nhZVb+euGCDbU5P6d2qQ2ixbUfi7qmQcxgFmDsFJYJc2ZgRJ3D5FZJO2q5ysb/nRm8Pg2dwV6xqH
w/LpmQFxckTU2fVqLW5Iw3wE1+RTdc8nYU/Z2PUwk58HxVyHSSa8u6tXsFMlxwbt9IP8jW5Z+2ZW
ycjq9C16f929QfYQPL5v6sdLb+MH8siaplB/EYMkOrcvAkIH8DXwWh2Gzd0/xOQ2Sknvk9BAa+fc
dSkP/RPMdyCiG9EEscXICzABpIDNVDFJq2rnGse74n2z4NHJarl4TSjxTJkXFV2qWPjvZn7Vm6Y4
eGNzr5XI2k6LxKGJDQumWb0FpEg/XXhNI7+dfMCQ7niLvK4LpVABO3sUp8nLYSO0IojFmGtVpG+G
goKNP/pFM6/0jfYgLZI2fBQApfT4libd0144bEwj6JGR4v1n4t3Pjmp6k8P2vzBc9NeIY6hZAMju
aHLiSk3IWDfndEa5GvXcnrEG8u8rkXMnW8vIbieTPU9ebqP0gY3ULJRoaaksqtv3Dbug4WPN0M4p
33aKgcZNGCof7Ohq8KE+JPVT3t6ZWJNETYtH9OOnu06Lx5JnblJOKmeBZkl3ZNwiAQdAVH/vDcy6
cASD4SeoXETByqdXVo/ItVQaqAlSYwS6rmaGAxyYDqV88fhrqFAthcUKKcbY1BPMRlC2iIBEt43v
yKX7fKxeWJyAaIln0p/RVS9ZP4Zo7zI9jBKzK434z5Oy0dEwSIo9KSUD1C4BRsJpJ4Lukxirwcm2
GbwRc/T2xaF6haWXawCXlKUAQ1RqDwedu7ij/FVpmLEtqYAgQpz5HzfzsgQnZMdAsy0AbGVKKmxv
VTm1I4oYldBsXRryfORXUwfvr94qYO6yqboEuqw1k6vzni526D6bf7Sal13g2y9Q9Yr6lfn1XjeQ
qRmbuW6sWFny5klAL4SZaPYHWf8IOeve7/dAZhsRVBikCVUx+FTfBfKk2zD2ptmXbFgkgbUaSPsF
nNpzWDaZoDGw8hqMA96z72fzj+mMqb+7u/rnFOiJwY5QyL/pTq4lxwQ1BS4U7M+X8lqtUYaw8+Iy
ubY2RsXO8viNIi10e5ujTyyCZ1f5j3vqKxP+3qAnHzgqY+OT4B3Vm5+gIg+2lM1CJgn9+fCLbcOt
JuoLOhMcU0ojhWfPGTb7Vu7LjqdNlWnRP7CQ3lOl2xyaK97sEUa5dk3quKSouv5uQpr4L7RTAVBA
2MdEpyjGiLvxYDH5MH5/R0Ynw+SK+/Zgq+/Qb6AmOz7xeiy4nj7l5lgkRtECEyFOwkJx8U0jInK2
YblaiTl7a+WuXYjCc2tEI62dVg9O312tSqn4ASo9dNutrIm3Xi9vGoPxKahSqiSAqBBMXbJQ6AT5
SIVX0Xc4fAH9UgCUwlVSB/cA4Sj4YFb/TvuExDcUPPNHUPRmFqa0md1RjqWH8IjPaWRYvzGi3WTK
T30WnNnhup8XE3PX8eiLNoojiMnZwHPnKdiz/o90ZIZ4rtvOBocP76kHMLqM66sI1bVE33BpTmBU
VB+gMkoKwU5hDocYaKENSrtp2uoc+bYfmFCx4wSn9aSR0MkSur59PvTAwmFGE8dK2/7n0VppJrub
SKtuAd9z0MuTAgWWcXDw/P2wJ+822UeoH2+xZGIglevtRDfbHVJe6f5hD+nmkYoDuVXJRut/yD6L
GyTeP4rH/YeOL+6FaX0dmYVzTTSZNZfMTkgNBDFnkdW8zdE4X1ZIkNVExMk47xNqR88tmtXzqSVh
nEsqd9uYiM6CeA9XCsRasQJwCsFZbNYDq1+mrk7Rtgjn/DbJJhZ4314vlYdo+wZoU2TJ8ZLg2Gyg
c6YCO83t7CoQ9l/0h9cIap7jxkPszQLHhKHn3Y+n3VcR8VkJKO+DL2MjnU0LFTyI1wG00RPQmfi1
6nlcQU1TzaYRMASAs7B+sq5m+T3ucVsbdekDJhPYlWrJGZGVyQN1FJkEbefE1dzupPQSN0AOVZG/
ANVcWV86wXob3xuBM2mhF0IvLM3rBr3HaXHpOa1Eih+drMdHj9mLSkiPby4ndpmBVLe2AgWRMoOO
6ddUoCOEn1QSHwdFxSEyrEK8Dsj7uFaeRRoFkQHiQx6iLcL87c719WRd764ZHOoNqMrCp7pZgd76
FL08dVCEQPF0GvY/u35Jf8SYfZAPB/src4lbQCPo2nFweCturKMWobryJrc/FCZqVU8s6wPBjSII
F9+FbLz6bmZGFUdVJfX7W80P4z2SxmoYRJ1/KQseX0OLS08CFURdJGU0VMvFELsVw7E5N4u7grpk
xi/bOP6tjl2enUao+EbXiuve2WBKrfZrhcGINfW3LJ5Q/cqlRDqw6JuJQFAjeGNqKmhsSOH8Va4p
yGCBcfqv9VpyxCV3hVPW69ue/V3pzHVwTm1CuRXX/0r5GyksK9pLAtwDO1/zusdZscm6A0gBlnde
3KaZ8lTJkDTCd4pXFSQBjsL88gDT2K+zRLGvWsVUvlEqSNTqQpPVCONfFfZNF5X5cl6c/w7/DrXg
Xf9u4b7NUn95Rk0U1hcUxoF8dOWD6Dj4dqKSG+PU8r7tTubbD79BgYjD0Zvx6IDmIXT4t142tzHh
8SguybEDVZQh5U8LxKiXiCKjCV+n2T3jJugK14p6RlXiJ1Fmlg0v23bVzG5iHWcKD+xmIzidqM0e
WGWN4WGds0jERKuGkI8gp685uuxngWvSurY7+ruR7MN6N7Co10goyHLm84dVSkBdok8r+pURVpUt
0vJk23MN4rBdBbwgRyiQHTiVDB98GeIoPPxEVYbPNod+F2MyrWDKpCgvoZwForcd+GJ/bNX426Lj
NUHVa0szh3UkjbwPAclYfXT8Fr69Yz0QUDlguuRhVWJymY1UZGxs98AyWwSDjOjQz7iRxcSE8SBS
9cIf1KlcVQmcoR66kWTV01fHmmsidQwznwaDM9Rhdg6z8myZrXlJUr1IVjc0N4QvCY8txHfBo/j7
ycXqnNbWHzMQlwLiKj53oitmoNRO0vQtG5qxfVrU5TdTJUx1pTdZPrVIkW5RSTqTp6aF+r1LwBuh
EwtcLWnVbdcYXhVuZ0wKS4j8BIeJ9gbd+c7JGt/7pkKUIKtn17Deuv5SeFn9EcpJWjG/N7MKwlkR
g3OpNvSkA97JW7MtnFP6Xue4phsGukK75Gw5WbOft7leyNgx9U+Mprw7Q0+r7HixuT1u0kZbX5n2
Z6k2i0yNgQ5M03a3bZYpTp/FCulgyKLF8f88sHeQa66LB/lxY6z0D/yco2qx3agYO7PjqBVqTw0T
NOtOOVg1RcV9gSnFSb8t/wWRZTR1qIOM2Ji2GAKgRfMdCYl7U0SmrDvq7+kk6+ZsgGhVQNJ+i2V7
H20FBLXFD7AiX8IytaXGAEu8haahVnxL1mNjd62CW8yh6DsYTz2t1/JQj/vM58X7O2SOVWpTmVIY
WnGDaHdyrUjxd9xaW+nd05fLlPwHYQiEmxEgEMWQm5NolLEQ0UbOT/1PAViyMhQXDPMcTAr+RurQ
g7jBBf0aoSJdErwKLAZzUkkjJ5zRpHHFIUO2bxPe1vCitYfPgaw5VQNp0oNWy6hQJgczneEvOcER
gC20cGOskYNQE3+/NceS8ADMZKg7di3bOe1F2L2UkLXZySy2QZjLi2SzV6ScbdMTBf+pxzUz2SCm
FqKycxtHyUyO1ntjI+cFykOi8xqLthGTnz1y3ot6SfQ8cnN9ga7wK3fzTmHk70NiYAfZHOeCC34/
MDr91S6MCudGOQMvPTSHFAAVwAtfGLONIA5JmVJ7GQeTXON9poARa5rhjNLpJF0O1t5gS6+bt8Hu
V3cvcLkOvmlgI0ePe2PR1KrUGB+uuq2HninItxNk4xmkin6kQZf+NzUvl/YepkN1b54FiOl3v3Dd
pZjKm/luU+2e9JWr3SdW5+KdtTjACY1rkuTVYn5u5V3/o7vAPnT1AZoy1dcfemdTPOe85BMvVPQr
tzV/TyzKYb+1D2mlsxasxjZLkiAa4kamaMiU1Y/KayPRYM+4IhkUdzQWiNSvJCllTm/n8Q+NF85O
kB6d7/LEGdNXdSjWc/NTQfbg1f+E3IKfJnJ2ReITPi940Gyv0TJh8O835ievhaf+HUn3oxvELBWm
fir+ynP31YITFmYg20RuGugTdCXX4Y1Xw8sHLolSjUs2KCOHp0W9tJaBKzs3OxZ9C48nYBrHQZmt
PZr0bcaWM3mhN/G5Q+WEQfAug69S9WZXzA8dZVn2GvZ76VBUAMelwBPUQHVhFOY/4LEp+uiNzkWc
92qtFhEErX/TgC1737DX8kLCG0M5spyv3G68TeUVtn7HlyhKjFQBex0QDJTwj4yRS7c1nEOyy9Zq
ymHmwfIcNZ4Xp433eXfdxUjwmxQ3P+MrIt+nHGgiY9KctNCqFPiRHdfIt744sT+l4+n2Mzs34p9i
sMjFh9lF79pwbqm1pjdj6uXyl3hxFnPaBxpmT9vse/yjR+bZHYzcJ7SiGyf0IPEe90QyWz6XbE2k
INdZGcMpRuMAS4lhFjKjhf9flQuGaC2mfenTFEC5niDwloUpUg1ECedCrK1Jq5wlVkHPsIYp1KkE
fWe0540W8LCdiU3D0F8bjqYtYVDqO1Ru9u/lM4A42ENnRIKda7T20d0KI6EWt3SKqsNw32vu40UC
qyYKhhk0XLhm0Fm0F8yRUWyrMRBtJyDoMbWqpvUUzLeJBr88iVF3hQrSBOzirLfe5GPqawRzHDPL
Cg7wQBKW7bipAR8lMQWqdhGpF56zASSaPtUfUtdOdoGNvaLiQbmMbKij2ZQMFfD0Uq2E8DxVM+KS
HitecSi1hfeoeqqP/awlfVEGiMG0QofVUDE9rY/mUmNkHJG37VBijIxemqFvUlbE+pPIxYw7LnqC
dU9SqpZBjFZLjbC5c6LjGrXo6jXRXOGKY20DGtkjuOuHGGQB3FrwEQYuSvzCKNBeInE2ypPMOObI
h4bhecw1amnQrRurU5VQ5ATyhd78/azT8FZvevHtXU0denJT3ud6laZTIBipuYIKFTFRZqhiO65w
Z86BST3UPPTaR8mLaaCDmvZCoUXkgzpA6p5mVsCxnnOkW/xo1dMmR4H4kb40Mh8rJqQHkiF05jWX
BGcnikcBzBrbS+d1hbM7Y9K6XDF5m8QmaRgrZrQLMvQxSlyMWr3PX8o7YpzVjkAD6zyllg+RC0mp
kfUfnfL/0MGxjgHDKrVlATuu2gT1naGSjWEG4nv43QhNpfjVMydiQm3fjIvOZFYUEMR4JhKcCU7a
7wW0q0JLCyJ75QQ7JcWZavhq2QhBa4l9qvFsf6hkn0GXrZcGv+H0AerPVBNcp2KApTK8Po190idm
jtqU43cfE1sz3wYpPrmvrU3xkMN5HjpXbtcIRpHarydpaQjJdsbLB5yaGRPI4C31MFeTt/39SD6c
0C4U0evF5dVAhBPVKOa/x+pywbGy0VHwW2YUm9AqQnXlS1LVKgJFoIOD1HndLpx/FJzuxV2MDSB8
DDdnjE+JsrNdMu2BT/9iNavB3u8gnqBHRHVaOE9FcmY0SZVuXiMy4Fa/LupsLJGQnQ3z5fYcjkzn
D7R6scX4dcTRChlitEsmN/GxXEtXeBJ1l1FmE0RtfgtiV5qrtKhVRiLqK628Ybj2cr1s2RUPYk73
v91zwux5wKPyLcRT/OI8kAiPmorWhkoUuEudA06iBGAKYISD67lQfjKPyviQ7w9qg2GmxOGseK8P
bstokynd0VQpTOm96A9qK3heAa1KnSM8tJaZ2Y7JRHKTpaBxg4pkztwmInYWEWj8DqkwPsa7nInV
NC4IHS6UfX91e9yF20gCV1ZrlSOS7SmcnRz+UAO9iwIyAhtj2EHNuHsUUw4WfjCxXOsamM0y8XqG
JNAUgKXbXwlhAG75uvilWN+WXy0Jafdkk2QfEAxFJ3KXjg122Qtbv9wCRqAnHjDKEAecQI1qwph1
u2D5DLR0pDzsKVSY6B+LObVUaIoM/jwnj/auIXxF921VgPjKGroF9TB4DTb0VMANTbIcWFNIfGBy
q2byXM1I2dn354n7e0Ow3BK2SOWPNlCJD5aKp0j4V/d4+tExBNY8a9TwMYIflsNBXVWBy5D787WJ
OjPe4zo+ExGqTClR7ov2Rbf36xB1t+xZkewSzhXtCzh9woNgUqaoYMcYFJTN2Kl1GiZtt+vKwE9M
gsSjjrFTtZjeVSRA5ooq4+Ny+ms1tscnwM6mk770yTFM7hMPSWT/KogxvPofDoWWbNimC0dNeDXU
XYJx1IdXmdqJSDTkX1sJyAUHHSAE2LHg9z9cF8jFwj4efKVvv5w0Ljl9k4QJNZQw7YozTyPA4ses
+giDAUGhGXxk4cOzyxrO9GcFDBzTa9tzHeTiWYM1+x2bPcaf4J0hQ5C2sxqfjCogZ1ZL0zoGm5tR
8ZjeZLp/NY0mE+4pMec5LE8gs5BtuxJLENT5p2mXigCL97fa8sD7lAqdCEyV3KLp9W1CMr++tJ8s
xLipc3ih5dd61dCRw4r0l8ykN1bGcVpuM0Z5GvJpDqM+r1wfSTBMHAdUUrh+Uk9ZPKjdPBQWlNa9
vmHdCYnc3PI1GQYRzuO4crG2d50HMsG/7PWxC25jQCnuz/1MnT7hrgVfFCqo/PNf31r4S7BwAlvh
F0LLkr0ypTflfwhII1mQO9hpj1Z9Yo6VJhf43eHsKSO0n3Vj2m0bvJlAydurWN8RCiODYP0OZ//V
tNt3VajA1wGgyoo6ahoj8OFE1TuefgT9jBNCdVlNJR2EbvjsQRTcaEtCyI5AY6epUUaZEVDHGwL6
dR6L9Lw4gyduRSc6XQoCvtTVXQyWOK4KabMpUW2imFn7PoTZxGikvicORa1ZgXDvKkCg9UD917L7
aWdoD+Y97gENUdqAcOM4kCynoJxGuFatoteW7dfLGNyIY6FSwsEiyzEEmsBcoFDR60WTiMLVGlga
LzALSuuzZFUEPkQN1zjac19CCEDubZ/5Xpmkp8MGFbhXert1CLI11AhuZCQWSmK1NRPJvsG7PmB6
2bVxygz4Jj7b5qFAIFhRP1CTu0falygQ/lUC44l95RzqmDwpjOO5e3nz04upEjyZPaeiAwC5zJnn
/oh/zrJ8EV18EQ86ttnWekjlyKjE2QS5V6qr53N7WAfgIbKZT5JI1aoK8trKJaOKae/+FmIREOgO
4RJce80JA8kIjN20P9uCMRpTlgtuRNGo7ipuv9Ii7N8AiJXWqhuFdqohM30vaYvZiT2mjUJMbhJQ
N8IFiw19oh5o8qm+KONN/46SAKvf7werzMwMduWyPVzBYFC8eCThEZhrXSBRrHfOpqoQ3paZTGyz
U2hUgATMCtEDHINPfp0gZny9HZI3bcwFBRRA0k9Dz/9jJdiS7GBFj3cH54xJ2JYPJlzJ/jUJU9Qm
uJfasIEWx9ehHpGeGfPnAkI/cus8nbTgvRS9p2rVvHbJeHmgFq6hp+Nv0kUTJbBJvx0SWXwU529p
4YLamdeeiTRH5jerZpN5j29hwBvZoVX7KJSMw/2NbdTAhygni7J8B+++un7Sx5cuh1G38GN+AaHa
BRDvvSXN6fzoO5wxOq4E8DG69odQ6WNdHkm7fB5QSF6f9vLQd3YMTGIgQSkF8wSGNq1A+7C6MSwt
4InbqupsMDZU4GZeMjE/aUXajQpDxA5de8EfPbd9ct3HB2YNDpo7tqFIHI1w74bVq1Drt+A46OeY
4QZIUEPsUkaBoaXTdOnNjTtCFgxwzTPeQhHrR0lCrSFDs9PVlII/TTqYtghT7GREbKcfbWwwVUe3
OuI+6AWEU04A/sGY+t2E/mVwNwp/RIg5oepGiLDDsIl77lwOmcJlO86Zsdkx4wOP5D0DaXtqWvlB
5F16pkVcsJgGvK/Vb7SIHYCWVG4ifdqcL0clcll/DF3/7Up/HM3jeXLH3o1Nfx6VW3CegMrOh9SL
611A3YWlz+FZyNp8t34ktYbA5O3j1HqgoKZR+qC35no42K65Pht3+XVwxYTnEjryF8Y98hpakqyT
LMnzP/GKhmXlyj9cnknL4lvymdeaFbZci3PIRPxReeyGtdBFHqJf5A9LLVGIckrFDkx7YkEmrFOU
anysExw2vh5f/Jzj43uXsmh4Swnf/xgj7dbO3UlAQv1puvNFWMW7UOmQF07h4gHglesuJPyLNoHh
PW+e3xNYBmcW808lXcj0gc3xnZPEhezajD4mgD4udo/Teyi2SVL/Pm1orkp9FcJt6ue4+hpFwsAU
yjoWzADuyivuC1Sf1OX5nP2yj3PHbbYM5snHjZPaSg+/gt+wqI5O4FxE4+w+9hLzlOJS4rI3HzJg
R93KRwJAnaI7LfQrwQVfTQ6/FXsL37B3udbC6DYKv7lIJZ705GLrnpiNmzcmXIqyBQ6ruS9ssddo
cCVjiYIXrV53CaqD3bKopdGTtYZnUJVF4m9yDPpeUDt78awIulQL4RqxaOpG441QWNT+sXL6+9v9
VCsa5LjhNpgp1Mwj1cv6Nx3HDIV0Ah0wOrkSHlHIL0IUQ0Y5qKDwdIkXAaHgkp9E2/1o2UmP58dY
D5Eh1rxuvRfU8ebuywmjLmTFjmTImqc4+uV4NLEnwhru+aKzzxa1Olbze2dY1iv/Htsxt60ldU+N
1icsgKaWSadeePxaS0EkQ2SbyCt0HKOx5xSYb2lI0iskyRXW3JRfBIBhrxbLna5bvvwCTTWGyg33
hT1HYl9ZcaP/TE+xDlKdSOYrQ8jIQAWrRCSLn2NoE7JzXqlZuXZEtFAPy/37KWWw6g3T1IF20iCn
H0rJmI6lfFqkz33fXsUFi8OBR02RtSWIL5rO+TCiK2DJjRv0oQ9z3LCUz6xe3BhDn6N3yKp3LZHT
6SPbGqhWLVWVbIvr0Rp8mMVyYsU6LrOBD7EpPEh6rpFc2tflHlZ+wZuLyIdv47Y5kyjsaNj9IKNp
2rQYQ1NvkwJFYXm7zfGquam4eOID4nrZm3Gq2GXWZyL4S9S4D7SdKH1E+FL76afi9pCTf4lygt+N
nmlSov6KeeH7zupYDDUkWp97Sv/MxZgEwm7vy48Kr5vNLf2CSQLg1DHy2WJDeB7wSa3sFWIHrzp1
hbjfKrhD1MgNU0TnW1xPSgZpe3RtKFkpQvoGsImmqD0rQ7oqvt+bFHMUp3acxKN2f6pdA9KbXVjK
7thszkwAPDoI0TI8gWprvvGify8PsT5uR2W9RVoDCmh0YJD/RH4lThmZrHLbu11/ar1PK/AtiEsI
jbI8p/N8Jp590mlHfJavZncQ3t9+OChe1pGvzJkPN7V2R8CnpEHCw7YEFDsMF9GRE6QeQmDQk8y6
+PsRWMGQFrDwpTnvupBJhlV0Dxd/LEOsbtmtbvS4a86nwHet8JnttnrFVXYD/zC6ozCmA7fP0qkI
3rGd9c9Jc9veQEJ5X0TpGEKaejAeOSjxOrM6S33njD7uO7zPwC60oslj+dfeWMqzH+hwtrRMeesL
weP+ZXWuLFcg5D0L+s2ORjRwYCxvlI0sGADzWaH8j/RCB3BjzYrEv1OtYV35+PYcKyQnlfROcf6+
zoeru1682efYcBYdSBe5cv8Am11Rt/3yXubaV+DMAlWlREAX4wNDBybnmaItyedGJUja5OyUFcDy
S/3s2d3bTQcGrjnfa5Hs+GEuEjJXCU1/v6iG8oVjJ9OED/g7JBp5I9/4X40iFOd2yGlg+Of9Gl21
EMi2079DfMx/hy4Px/l5pOp1C6+CP4KD/Ifc/L/tRRRlqV6oBnGGkoLKsHQt6qHK2pvkNfQFh6BA
N0kU7QnBYzVpaBsgvbMt2o/VHJQBPmDAWsanlHR9m6YruNk5Y5I9K9gyQ5sLrFK1PJvqGq+reJ99
zkUhJWYsIK6RcWst6MSzo/Izjj8vwZp7HQjCdO0linK8v+l/ndQwdhdpy2UOYGag1nWuwmwwMjrU
Ne5UKp10KvjFpP+h4wgQhR4WQygEhG2Uz7FfRHrTTIA8IgSRBmNDKDW5ii+yP46GInNpGw4ZMkRv
33GPkNPlQ8leuzZMU3rvZGmry8sef8hHhHCH4AdfzJkAoU0QqpDzka+5k3cagm0C3geyK6zzKZ4/
d+bVPELJse+YcmUgtPzNRn3g3obzA8eIUTn74L815YQHp6WVufrE0N5DdKPqjt5inD3dyMPFtlgo
L9dmO0B2SFvAZEbJ+b8lhuAls0DLTtw1HiistFpSNaXa5Czk/QH3Z77WR8l8EjqeM3/KXhK4kcMD
yrVIas2ytek0BJ2RQKMyzjOEj0O8DesVg0QxlDg1NMBjlcLoXwt4BHYy0u4j4BN+1j2Gufls0YUw
y3D9E0dAU6ew3+Qi2sU3lggsxNeEylPYzShVTjgZTvUoBPA6ePJGHFmb7Rzgrjx9e9CXcMR36vMY
kvxhV3XM00OBp/PfdwzXEVA/Mt8PheWVafIH8UWJtUPfLtEtokaPlI0R4NbxKwnYfG2KXwF1uSJR
zBKaunhyr5vj2vGn2F9muTfMhCBuRviS2TF78FP6cQong8zGiNLBNtQAkYIM+fbCqAmORnjtlUUd
b1y+DObjlCuhW7q6oeftRiuh1ZJXWm6Lhj1KFbguYodqasl/W+nUUtYpYu9x+5QWekyNSbqGD8Ly
O7yVNwdDi8bVvFnSk5WaiDXp9xG64LGKd5lxykE1e4MTPd1uLTVxqRqypotLkzchZLSVxJp+6Dn/
kQSYZ1c5DOuFc3sFG3Fpf7DIHrpYt0mIczmEIWA1sAwMnsNm/wFTphuh15uckhA1ImXSiQJxFTaa
cO5fMDSQf2IkEju4VQQpzuQKAZlMSspjNcXSLDb6z97m6bcOlnNZj63hIFcXuu9Aw+JA8yYIb8FO
0IHdruE7GfyfiPCu8NFWliCZcftxxwSYH2DjqHV8PSbRPuwxTawJSYI6KqM/cJf7xHjkhquqCAm1
v+/UkwcNbicZnOa8rk5/PQxZCBf9hkDuj9/2xrFhsny+AWalzi6TRmRTJnrEzjgIP/eyW6ItfNaF
jbnjunHJEmx013J2qdXR6MCPLGNOsHOGXfbH9LXO+RBj7IB5E1xbmS8KcwBlD4r/fQRfdCIAuxyM
bMTzEe5FD9H5xtHfpsuKK1ATWa5da88aqoO4IvQUpjkZ1bxpWwgUovQwO2NcaIwhTYjA6uApSaiQ
pLl8Y1nyNXHS+lSLcMAD6NrbyhSAWId2mVzkqzbDC2ELXB45ZFt3S6+kdXXm3fUhFc3slY4Tg1fs
SDPUr28tRz0yEMkL5aYv4+FOTPxqyd3EFIDVK56MI5gukzNGhNBjKZhG7QSdRGI3j9NwRFyRcnNl
9nH3X4uoWcXYMkh1mKcb8wqO8WAOuogoe2dOg+AYGBVbTZRUhJjMN39+TXYtVXwEc9TxxYyJoGnt
3x0S2x78trh/rept6w4IkTxS/gpIQTw4xc1MQewoLgZrk5yX3zmLZDnDxFpCkrmAs7xM+24NW7yU
DNWSBEeGyHvbd+ThTytmV17yrqVxk2eVAiKBF0dVU2d81vkZUNzjiSOhsI6m5lfRz2qdMfwWnKCG
hqgxQwZulu5e1XIvvHokbzJKZxU+HPG2SpsaoATr7CliKdV1XsT7YVf7uvRP9HjRC1Xgz8gCJ3G3
ib5DAOQgyAq4OrnQyjCCR30kRHgBA2EHMUuYSdpEd6uqZkAMqRNcdmplCkvwWju7MBJz7SjTObZK
p5ARiqgjMj3HxbG3950P1VFTo5DpQSh2BQez6ADDjMe64097Pp2DxzFepX84uqj1ELWmRQiaqxH+
mvDYtbeDXCvy4Jqq/olJ4ePSQxwRa2Vuet8BOr02jwLj8t99gzBzO23TnRB0XfU+LbsP699hfsik
CbvZwOC42PSGpic1lRcrk71YpCb2dda5yEJq9IPxjVrwaywKyOq+RXoIzogNp8QYWYe3d4VgxmSP
cCptj73xrzuPtcIVTEztn9WYLO8+tdQAesRA3ydIohjyWdOlAqh+NJb3XnpbncZ6NRumHxz7dDhM
LyLUqA4siMPPvuV4GvCPDssdwWVZS5C6cFDEPAQQ7SMPtJGttp14/wnFAWeMqKWwk0WSgjoXgrrF
W0BPaq2dCZkYEcs01RqCMXEUdPGkonSwSmd06gaoUCrFsWNd39XoC9k55yMg/2gOvZK8Bx289hQN
wDBdpy0fEkIFT1ZXNtM/PGIvY6/yEc00Wu2kxsNTaCZ+b9tksSUrjT1h2idk0a4U17HSObnOFeWp
jn6kMw9B6Oy2Cc1pmubZ5pJhi4RGt2vHOuGgLB+c5euUd4I/U1TqBKf8L1pLoiQfkgD/A1slcnAG
W7+GcGZihb6VGsvaDBpuyjFaQ1s8EDLauW+1Cf0AGT+HGLzDtEaCOx7FIS3Gjr6O/E7Xa0Pgv8zm
18Jzmnqr7nbtyHLVthQ0kZfKpWIAuZWJtpePupLQh6JZi0a5gyafd9c+FwsjKhQubJpvQc5ZyYAG
0kZ6iDUFLMLbZktjaJiJ3qQrDCYGEYGA+78XnMZJW2na7ohkPQAbc1/tQwP8ON1wGmQ/IGv1FFyh
rE5PyCSYvjEQnlRgCh/QYxf1bM57Z+sGme+RFXxWkI0exmQQ9UGeNgbRkjk1utbJCMKBd17Dig2s
KNZuS+91oK6tq07EOYqZ6PVGhcwqshf9YiFM+2BEggjbyLMbRGp9Cp8H8GEanqxIM8rro0e6kUG6
gYzDH0W4Lk4dIk0A+PCF9iev1kQPpN8WlQJuDnk06iz9ozj/Z8ozHC/mwuBNEpngMPZ5xoSCoyrb
2lzA9nv/rxE/z2vo9ZGgWdlp1RdY4by4id8I+E6k7vPRE2FnvqewH3LncbexkjcAZ5zMPu+l3G0L
aymBWy/qzXF7NKip+4arD519W8JSNwGGmNBYknzN/2acUfKRs7xw6Y1YkG+nJb73+UpoOr7rFG6N
6Pk4YuJvhW3nA3r6+5AtRbwDEpmRByC1LaDWKCSZ9I+Frqi4hZVGbFf50Lb5eO47RCQ0uKd66LCZ
SjImyo+8Kv7/vf3rCHSSu9sYuP9445JDYwtRlsMhiCBf5642TvLXZSY4STyDOBT/09h8nVWLdfFz
y0QOWOiMrbQF4wSq+FXv872tfP87fHgUTf0/mGGb9nBt2E9xYBPVfy5BZibLV+0KCkERynadydb3
jW9FgO2JRJ+9qAqfQH3ZXRP+NVmZTT99wZgbj8bMgu7mRZhPlgU6Xt5doBLTe6YVs37jgQe3ZIFg
oLCggtNWgJW9grE5UIunxiWUYD4Ne3cuIJv+uOx/Sxf09p7e8Urgo7+dUVxdVqndq4lJbfOHATLc
9pDByklKX9Bn1+dJtid3QtzhNNG0jWScN6B8ndmWTOyUs262C7yjhEwMKNJIetrGyrg0YcnXiqYF
AfoikcFJGLocY5Ux/mcicDN31Ixu15OSj7MEodNCXGMsRhPt38M55Xs36J5kziSFzwWPIQ2tqS9u
hnSGhd1W8cOvoYDTrXTZQvyYFH52kjp3fIgkjgbJz6ajgNS29tOENin5971vBk2SQdUxK1vVqcZF
WuYk8GRteIn2taZ7BSUO3SE7kvESzdAc6dFkFtLkODXqavj1Tk1uB+NfagXG22FfbcHq57iKFDTg
xUO45N5ZMjhLxjVUZtdSxmMt+6S4QWP3Kgu6U1PJC/SQKiPApzTkcKxOxM7+/cBaw1D+rxbG3vsC
UA5pxweb2VjG/EzINNWPYHOyqRNYp3DFHIOYDlnIL5HrswG0/o0TGiweQONwxRujEkIF6mijpUNw
rsAG+T1KQqWSY4RtjQuD1NX51HepkY35CeiFDQaX732jm7K5mb5087mhW2fQEhncvQvY2sq4X8aJ
ZBUi2mPsI14PnGeHmyTU2nM0o6y92sBxgTUVz4UaFWXadFn/kvOIbqEEwrgNMvDN1hr15lzt6rVD
UCc6OAejWqB49xNo030z6oR6tzLtGPBF0akhsb3IrYb7abO3nLLO50cQZ7ZhW7jT9AuLpdD86tKV
HPcLO6WiuK/UF+3N7iF/uWtpDBnQHv23EK9dfQ6pxV0Qg41ZFdNLFDf4wY633NCxAx8F5HY6WG30
4kRiB47EY1qDsBrnhq8/7TSSe+C+Hf0AcjQ49dc/5pFhetaGbHi9f3dFKCssSir9QCbI9z4yr4pd
+SaizPyZj+oBVt2CcGyo4OvA72dHCHhqdz7IzyBwnnWil8iIdOkBwM39+21PXXgcynYlXxjlpmNc
6Mhuz9M8evpEHXKoG2IX2WvI25P6nsfWXMm+rYsRzFO+Gvu7tRf3CRknC9uGailSgbOxXV4wgkLV
owZDqmHET5/e0/Dh0wsWp96zOEpUxHh21WZtTVgZmktwL/B+8xh8PC0C7HXDVzrPHh3H467jfnT6
Q8NbHM+4CnE41WdhYE/PzCxBvLyqtG5ZQpfFmIMUqK5iButirl1rjSwa/0EeYd8hcaBJurjVZLhb
pIOPG0VfOrwJI4qLpCMvJqUgNBqRJyzoCXL84w13/92MbUksq7jJ8NWIQ3Y2YuBYHzWqYT3eD+9d
mE/1BicYj/nEeNWjwCEmjog4OR6MYfyLitrT83RKmYXWADQgjr0/5RiZH6mr3Tn+jHcxb7bEus5e
ND9+4g6dSl1eS8wm4b4L5k+e0EDPKFcLcv4jmf6aSnzdo182zh1wQVS37te7jx+mJCpAUJGiwOAk
mbsZnoIJRsV01qTTez2fa1O6pJkrweTqrYB+I1dUE9Y90wRZNsHWN8mvyS/7bNsagLdzWQLLmGnV
KOtAB3VGgeikeM8UdOGxibOb2BGQajqMUFL2O8FiBkXNjwadeuUdlRhIA+LMihT8CzIXKHaHaQSo
XQ43W8RKFY6EC0ixkOD3F+fzbh6EPMx7FthrdVfKD98z6VJp/vNgA1KDVmoOg9OZsVBRKwCIiyNC
pAXyqemKCBs9kawCrokR2viwF4PjFBDl2LP1R2bv/+fBugR/74MQYoMIMihQg3r09YfPvZKIeObw
9HcREKzCsMKbc5yxE7J98zybjp/Kzl4Ten8aRLHSKuDRXGSiw8JdUtCmS/u81XXnC3+oKbHA57SQ
ak2J9kZaSE7xy1X4Fb4yI/qDtWn5sSx+ytdk5xLRdcER2u2hkCtekVWjsIWbcUQExyCPzJvVazBP
RNQ49+PiB0CqG9V8ENmUten50N+hkpvp2SOt8t133aSZS234XLu0ZCPm7brjVH47ujbxWez80ABD
C/DlhOahswvQBU4fmlsTB8dNlsc9W6kdmPdvaqHe67PfHlK9G27YR9zXlL+tdGro6RHYlWYz5iFw
2GMssrxuxG5tfKnT6tACdR17/O+mX7A03wYF0EK43d+7IWBgARxODAqSFb1Cb5++KNTfwMUQKY2o
mVr/lb2RgfUvAZU0gE73EE/yauAxrZAut9zVRpx2KEgA/Qc3MPTI6esl4aCLUIeqfAsBepuhL/L2
5hmtMXBqvtYbRNbxp6QZAGkv+N5BZZMA3nAgqEk9WdA8yqvyqHEAnaoQIcNv0q/c4WOoHIAU3xg0
zQQYhJDt5CaqwPg2eqRVyB7MHNHkxXDjOFW//i5LIeLJvBpyYglgZKtv8L5a1b97MwZJ5dC6c7FA
uQ777TStWmkUaj5pe+CtlvxzXLMVMWjzE2QEF8FY0rRZAkstd+Tgc0PhWQOTQjefS+LOQH5MvTbG
PcesejcdcFfQvuMqQSiGrEC8ePVjH4N8nxKDDqn9KOImwLRll4BqqNPSdkjiLGbBrQu/amUUFOe8
uQvtFC+OiXyJG0pDiFans0msNIAmiY4EESe/gWGlO4gKmX+/GJLvrx4Sy5NWCXNzFHrel2uJnhaB
AUI6G+ZxM3A6D2fSEItMnXshrmvJZIMuAt43LTC+BSLRPZB+m1gkTAHacr1XE9atZF7Vs+EuqPLi
LXiaW+Ck/njdfW1RvZrb/DcMSJSXJXcyjShH211lm3nuFHUhSdLd3v64oVoB9qVDdXT2Ct04o4y1
OP4/wG7OqzQFJMedw5IYz/8M/TFHXVZ3GQ4L+03ZFvHyxv7WqjHyfn4UxYbvIHHC47ygQOXyrKJy
nstX0L/e1txloOAyDng7pY3UeMRlcVdk5SKGrpqkdbW70CbbXmxwzoYfLbImaBl/w4vzCGP9hO+E
GdMGStuBpp9qo78ZsNqbk7FnrQt3m1mi65qmVht7zCzMCzz18gc22IsqMuyVTeLIZ7j+urqY2Ns4
cjPbZtutmXDP8DV0vhaPO1f0bEApNks8u6IJwg8jmKosdbou+0MYSLcDuJN5x5I4eUlRxRWYhZwM
W4WpSnuuv+Cv9aMy9TZ/FcORkMhi6g7Qvfq08dws5LsAN45LT8N8dHcCXN2Pfjzi7X1mS6vPgKLC
9xqRpWMEQcRgyV5TCmzxOZO/dPIgEhMqY0k4vSrqxiZ3F3eX0A2CvsnxGSw62NB2KzJX4owBACOi
VKNEbsZkQnL0LBvtKJidrTekb+6VseNzVcS13ayxXJTpv36lFiRZniIlNg1qf2f10qN+mgOWkcLR
99fLZnxpoXR6iDlvL5Mui67zyyKZF3VSMqhRm2HeWCZZATOEo/wopRwh7niNM4YBd780yKm5geWh
Ozf9kYJrxiOzxDiKMkK+JpWUC208hL3MKUD8eQmAao7dbboCBOJV3TUqJwJr7AYt574e3gW8QOa3
7rYuJCpiA5p5poOIlocWnl3wHuaz07OXwgs1eSp2zXv1UlvvC1DTmYoozNHVNGDb+Dg94vVbdKJV
2adyl0sto6GfQCOksf2xJanzYRrIScVDZK3eXVBawGx/rYVrgREIWBBwFQLwxCPp4ljGIo12kic3
gAqofvce62KdUn2qVKBxjK5xQgOwsR/Dv5O1wsH7loRRCdH+4eSQzpmemD0vCsjASIB4FPkdI3gH
DkKxRAD/jF92EOQqitZ+f28qQnux0tQTRNs+dk73XxJrhHZ3NCsAB0G7qrcPAJDYOn/sowLSB2Pn
CCBlJHBQygfVR9RDNVtp2Mknr9RN+GYKBhceuJQVG6H9eWwDmGiB+7rFEXXPdXfggsuaQlcvEvLd
Jp1r98btUQ8sG9Qhqp0eBSd5JR8YfMg6lQKfepqe0aXsAPzOzmVuGBDrzXbIqayK3TUm4xYl7cEJ
8qvVmHsaXSTn42aQijhEA342w6v/wkrc2mfCeKsk8NfltTBbnjMeBcPK3IwYuwnUbdh/QnbFTzqN
Y9Di5QsTrnkJ/n2m26QewjPUxFAl+wC5fji7yIjROYctTDJYPJNMPHNe8HdOUm3967BlGknpKFkL
oLp2vcC8P/KgG6F9IstYTnnGWG9BWYadAVYUq1pprNlH5jNBDR1vjaOWCbmUHsLiUoXSAARtmWhY
4D96aSdSUit1BNhHKrszaE/a+Rgvz6GHbSaPyuH6sR+hYpSTsfR+ZscBhQYXBchxroqPIvsEitkZ
s7KrBsmgPHw9gIKgD6H3NOQp1bcpUuzLedaapvIWGhsxIjWjtrq/TaxCQBpkBOO31fwYuMx3MrjX
hKPSYrnlF7OngQLN/W9ct48SbU+NnHro841HggiVSzA149QywJ2BXPb22lVAvVZoBB0rNt31GxTE
hG4Qu5hZnJoeQa6CpWlARKxWTfLLeA67pfW9sW01OFwqbxjiP92gJkuWCgq8myJwHKALB0/w4C4Q
MvkdA4B39rI/H4L1mi8djUWJv2ewcCL6rSkBgAxSwI/A08BuxaQaKFv+2LLwHrI2dx04AlsWRLwk
Ll7MdP8Dx7cJk0jmxwLTJoSmH/dsxsVCC78U0Z3zWffsTinDfFnJ12/pZYdPFhgO18nejfvQ6ax2
Oy0x65qYmAoyg7a20eNPjRXr8/y6UMymuuBhy18ij1nwcZksKi/8DHwBZMveyhRtBDFqrHdQdr7j
7lnV+oj0k27Yyt4zbWIqeXZHyfaCiSjo1+AyVZCjHJ9aFdbz+OLUeuLBQYJ5XSWaQP7kBRi6M+nv
Jvyn6QdN9FA+cjKE8ynTTQXIL52Fk3ZhakPJHcAeEGsBHovehKvH+KzeLNq+0RRtZ/FeP5y+WUiI
Yaistoyoycv4UguLTHt8vg3kxXREzR5h61YsVE2m9wW1w/p/53KCbOKrQoeAEbYLpysNjfaQd/Dc
oly449k7gVRoL9TZhLuhDjBrlp2ZOoh/R/Susw4h7BXcQFQY2qUXYZVFpkM5j3xs1yhn9gdIRuQq
5QZg4D/pR3ukFeIWRGFi/BYBzBlEAunZHtExGfTl6VFXE9LzoR/9PISdOOyYzSjTCfAiThA1OlqC
5+rl8NhRKPNQ/jHQiE5AJeCFQPlxs0enIhViglxRGvbs3T1FsHxhTcQMFQpHOodmS3WGRhb0BD0x
OwgYv4pGwWjQuCuIgg7agS3DjOUYjH7ApFrendilw8Sff76pBEk6ElYwZeC7QQu0pugYgvvoMi+E
K+IrpybT7XWarHqL1KOkm92++Fbx9rZ0FiLYBTdYz2/VHx+wynEvLzBRumlKGn1fjsJdWwQb6M8F
U1VTEVThD1MWulv/fiSGlxd6FjHwN1I2ewkhNlQg57pJyITEHa7Z4OvjKtJ79gdo7Agpv79B9KeD
bqkBwfdThJAhvsfEutRdDRT5uTR8L38OT9PJBXmNJc6TT6g7Y+v1/rgmDSPsrh2VIHuC/l01aq+b
gN0kxJ5G7mKb3F+lcvgnSv9DlvMwBMsSkr0cIc5qlxB1dachH4HxF6V3v/WhICA3wh42N7cBEqJE
sePsKY4qADiFFoMYUsgPRaFSKMWCDP5Nym2aaN1MCRgz1Bs2sWHAK+7hFkgFSpdL6oKAysLxiDQm
A0PAAEJk8zzMAc9ev0ZOaw0RqAP+7ZOfCG0Ce2rR2I/s1VUpMkch7k3z9GreSyRTV0T3hBD1uxBn
ZsEE/o/pLw3oILQziMr9YkKjoFvM0fc5eQyMP2UWK/MJaX50hSpkI42VVV+fym5ZgrVI0KlgfXPM
jXKrZEvDhAcveyMpyh1aNZGTwBpmMdXOCIohVag+0b4jGqtXFyC/OsnX1f7YZ0AvxPf03RNEdcUy
iRgpOXHoVDgSIMn0hDpDLuFYR2FCC9PIc41lAnTMaDtXR36DO30iHokjYRvaPfgyuzMNDiai4cag
/EdbhN0BzZhk2r8mj2Ojpdv2A/GQgZkmHFZYPdZEahsKtu1pZpTMA/oM+i2xFBS/Ci2RkqqO9sep
SyjFRDufcPjZj3T0eXWRcSfx0W0qoWL6gKGTdqVtjsCiEoyTIgWMKyN7pD1pWm5k3X5uW7t48eV3
Jiwix6ywTj0ed4g/ba7FzcaAOKmdeDXmKqcPAspocEIr7dDmUTfaCWvLBISB8YbEORVWRGOSXSyQ
nEahyF9OXJpjjq2ReF6jBzFT+om6GZ75qiCjKGCg/PxKaqdMDiii9MX3Q5vvqoA3MG+F9s75z2Rv
2kj34sRPTcbBBhsXkcAYTWx9kMGMiRPD/AyNGmv+K169aJ70+QJOX1/IjNStOvE8dTW63N/XcOUS
l3dIwYlRyXIw0ownPRnUzFgKx/XH6BKGmBS+FIuMFHYVBSAtHNae7N726XUv0RIsCv0XrLGLHUxd
fJUnGGbcQ4lelmMEFBgiXIj/V+rf2vk95WagxCWdWnaScIdorTHHKmbaAdpJAGNMGkhYieKWwtzP
y9AEjQsp+Csynnp6bgVcHd/hkIpYaSYRIi9NeARhIfa3b8tLvajvAQ+gH5SY1zOM0WX+S06EHcar
+8B2svwJp+WQ8YcEIRnuWv+IHm4dEORFONIIOFStwkxiFa/YmHfI12supixEHS0AsO0aGWZ7QeTB
Ma5RRurNZ79Zn/11w8V5iUanlmlD7hSmeOVGTi+P9LI4XK6uuJlk8SJz96HZl3qKdYx+11cLnuhP
osOrmS6vd1sw9QX+WNmsIEdNeN9dadKDOzweHMSEr+y7g0kmk+yBWlsLOMUZ1MNxAPyn/IC7JT74
/4wg8FcimqQSh8uRwd/VT41YC3s+j0qhAdjB9iIYfQlk5gy5g3tLXDX7HOrP6v2/lRsvmCbUFmpO
aISB+YcTuXjY7gVjG5r6vNUOrkaTY9U96HCqDl1uabE24wkySTXY6VcCGQKe42oAi46Yl1DPZ9aW
AR/lhZ66/U1eiFV0+osLfhXTjg88Nv/lkjqRd9O1lnV9fo9Q9dA1Jmd9SegiP6IrmNKQdmgsw97N
AS+aMoVoz1RrrVRQQVZm2x/bT4o9PkLtawdTNKOPIyFi0Ce/K2J5WO3+HB9Inptl/WttMisF0fOc
KTcKBHpKEijXwG3opUGicw49SiOuHWrUto1Y5l+uMWCFGwrkEnplu9zcXrbzCEBEqhNrgcnQh3Nd
jydCBtNARKo781siJovFWMKWHuEWd7ZNn83MJb1rOgQynDdMSyQgx/mNww/H8Igh2O6DqllWPujX
SU4QLhr44/eoV+elvSLGpGAhVl2ANBuqqkTbQmJkuBXcTLXBzgMAozWxcVq6rqqRkf0jBMMmHLXW
oWmHnnna5fCfQSM5hwwfFZFLxS5lPY1AunecPUAgbuKgwPEX0P7uPqN9Y3LTS4ZJpVKVXXsEake4
+ilCoD+MIRxN8dOHqbWRERkSOsqmZoAkGl5KpB3IKZ9qYok9tOhiXYrsqskq0ZwmUcYVh52PmyOo
IgZSmFnbIj6jDuVuHkL26rYui5uk00vRfmBKmnFaFu1rmMW55fcxIFbJpHbjpLOaX5WgyFDR0FRn
Q5EWqd7Nr0glHzyjUT4AwQcy2Y0EM87xu3vg8BwqrzS3Bg2i/TT3XV7trxfn32hM3ZPdUC95tn7X
64Swm6k7Sqa+1irpSmeH+YlK3r619SElmBXC8nt0p+yegiLyHug6Gn9VvfDhiKF31lhOOpV7AGaj
rG9DoTAYKVOZkSHMwjRkjjqYk6pM4SxYhrvbyQNQWXhy4D2T9SdD5R80dlUl/baQWQmU4+/SwGZL
MugFvDaJFAT9OMA1K/2pYZz2pECQFXT90aL+/7tGi8m2wtVdVQzcYXLQT7ZpWY8EPG8vowysY+zO
Ak5cucLGoDyBdW5sND/8whGdc0uXkPmFQAHDbUYlf+pmRl8MM+kAzWoHhfAbpJcH2X/yuuzYsbmM
Lyhn5CguFAgU1KCVMhzK41IdFQwQkjJNPtSJlwCQRZWKvKrQLFVox1bLqmygoiGeO6HdWYyT6UOF
9JrkkzpWDnEj/WtOCDvcCgFcgatw/qQiOdUVAg4Tpo+WRHeWhbRkB21lQYFUnY1jHyQIzbslkrEh
gKVlTA6kI7sGGheI4gzYyro6Zp8YhYm5AGwsbd9K7VGzsMI3zoFA6d9zcHVa+w74rFPxicbLAkJB
brLXFXFmIL8ccz8dQkpp6HfBBRDYd2rC/K1vXRyoK09H6v2gvQkHv3iBXUAmXG9xO/VG9ECdVikE
gd80LeepRFRKq4wnYajELGNq8pkYZhNVnCNLbSWlpNvVwZ63GQM9oSfKQQqjsIDRH1o+7s8wZ34O
tv6Gp1Q1tRnifuu5t/JuuACOceJSOal32XrnGJQ67qHyhy+34kdrY5APtuCu9ybZF5nNV/NWr6rA
Y+1TQuvEIaIhx4ihwB/vS6XqMqJ3NFHlysvtbsUJKlGYTQSWA0hcNCpPzEP4uGGVT08WO57Wtjha
BOL08aHovEbO9HePCx4bXmEgnt2SI62a8M2/pAoJ8G+5XEY0Nbak5tKQ1tKIk6Ihl4b+UPBwRmC3
s5lrZrDIsDJtDE2p+VvwO3pQ9ddW+hoTdqRImMmNyopVvFpczqnKMKLkd7JttpL20+ARmeHI8lKC
2SPlcWYDWNFKYEYt6QTPC8Tfqowqs0Si1Rqa50WzeXaI0Qlb9TJG/DCvopQ3TjrHKrg1nxAwt0kI
qIl4Jp877ENjMKHkQreMX3kUh/1AeNjyJwPJ0KwHqlnets01rCHaRbuMiyy3UADSZNzsoVG8BlYb
3Ddb/HBRe86+/5jGHw08q515G+dgGH0kYZ7mT94iaQb0rJ2SjCgqwv7WWXK74RcaRjiDIXIdzSnc
OztYdWT/ffjQWDHdow5oZ3H9fssNbfEuQNH8CsUjc8UAp5cYPYIFjeDzA1jWpDIEVCBCCuXLbibI
wDdNRILlTAPxbkUcJ6l3441hqRwu51coUz4h4LrxvNlFazVnEJC2YZ23AJrnjROYlEqrSyT22cT/
CmLqRS5tzxxizQLd1MxoDzlOo4C9jHvJ94V/5MNsMn1yIQF31JSpzst5TbQWIx8Z81GM9Xz0ySod
jOqbFi/Q+1ujysSqu4YGIo3ktjWGr6NIjk3Q1kldqym/z5zmNLUOucOwL9D5OLBR5/iNOvrOBvgA
gnij5MLwfar3aR1ilmyiI1LSafvfeX2g6dx3yb/3ryWDOrJjkW5kGOT0MZM2++X+RkqvbngAMCwN
sdNPBQ3xVNsIGnCxINfbYl/8hzeog5afPaoV0u9os8kE5V4FXv2ZWKZWGQ0gY3JfryYGoM/5LFZf
7AJuOnUPq9e9bBTYwSkojVFbD6sm0ghONbO42R9SwB9B2ZPG2DG00C7i0tx0KpwwXjABcSsFc/N8
N3SY54v1VueCY/k0WH5eFlCTWwu9FqhVhyheFe9ZltP3hj6xGsKnvLTkBDM+FDC+tJz6RS1oGiI6
+E40B6UTHyktctUVyKOIyf9VsWvafddalwDN+O1FsZ0Vuj0pBFP+faQ3UEApX6MRZvtnYAwTJvN4
AgXiLFhJomJaicUeWY757pW1JZR8VevAQsEayRq8vQwEn8wBhZl2SG8Fa6KUyA2HAaW/R2Wmcy9b
gbeGhdLP772QstA9fFcqvancFXhfNZMOIWN1xSW/GLSpGCgMFQIn631o5VwSrAp7YcDdTF4eQQ6H
FRwtY8yqfyoj6FX13jaDAQIKmeWT67nJ1qnzPx5U9G1aOkf4m0CBDPvuFpaaZ+HZNIGS2k2TLJTt
xp4+LiRGE8zRelxYNk6gumJrmx6MVnyNKlioCXVNYJg27ZzB5onk2eKa+Vv10MsnQ3g7RpzietQ0
6klupXq4F1t+VM9nPP2bAKRHcXbJzrgl+aIMuMpnrM0adwGF+97N+MFFyz52nlrzdpfoaDttBILa
5SZKg5svAqKqjNa9rS2yIfRVLaPe5d31EY8QXXeWBCimyW4ZthjvCwl+VGg4b5BfGTGO2L9uu9z2
sDdiC21smLHlHm9PH86/IA4vfWabXpzfV4KMd7HAGJUpTf31VkFjP9AH+ioXFPyFbiY28Z0x7WnZ
KCYVGp/RVGMkZAUcJl3VMamIoDeKG8miKav8kGTynuMrlUwL4zPR31eg0xmAZQXo+8VUZCKD/jTC
Izy+9bcs2dkZTkWoZbYBuoDjTvfP8j1gSm3qA88aoxrE0IC/tjY1ODcT7h8J6DCAkT89qx/JaMbK
uXfgZ1znHaA+Zn74CItUYki0j/UreuLrmmvAXvpMCnxgIg0hDj94/SuGYup1U8Pw2Bj2NveeH0I6
HGedQTT8HmVBeByyx3RpL+RD8Sr912YhBbqBXiQ/0jmIu6VsKILqq8noh6yj/E6vg7iOQ4yYR/QJ
Yfxz5OxpswcOZt7nDi0C6xZ1Rn7P9VkSqjAs31mkxeCYyIh/YTC2w4UDr/0BOwmxdjBXLDDeH4H3
Y9ZgCoIR1+RI/11uM7X8OCGwDwmUy+jiMbvqXkjMQF4bpTGaDDcPgG1dxjgRsMKVPny9YF2HdMyc
TQqGahwEq69oQ7wZeFhQEiLiATkN62BzQUvFmkYW8PZk9kO6R41eVKV5E9JCXm9cwpivDw2yo7y+
/qWgitNX0tQZmxYsQRfE2ug/lGIxyoAuhzYsqnOwZ9j9cAt4NjYOreKxLl8ds8OH/WoJ/oy/OvAi
0eFxYkKE/9V6x/qDqztqMqhm4t4a9JMaW60hU85v8mahKMyJWbH0Uwx2WPZMJGdaDMPOumAKTEPF
uKYyFTnL5bNVS4fOLs2w4ESKu5oKfw/uheOO1oB7pG6AYCIVkT2sTXtpmuZ6fzRD2yO89wzqVkO5
Q67KKIq+8fGiF0UdgpmXL0fwkZNdkxKNmts46886Af/KJNBxy06R5/Y20pIvGvup+TCylNWyLY4s
+6KO9i63LKT8AcQmUXXMzJRnjyzkKw/2NlL7gfAQoDF/cC40/Tvj6OS7wzLBxSW5LDBcwltihUsY
wu2tVrsymqwzSnwp93vZPDb0AaygPxONpZlMdg6Xv5r8f29YoiVI3ClSwMCgxFrui7Ah/d6UhNgS
mGsAvIILs/RiJzjjtCEf5qie/+iYdBBcttFRnAnovvCJjmn0KGcZ3AbnSgrA3GVbPnnRqTGbw5gz
P71w17MgLKTAA+/5nWovmDMyr6CDKrz3DWFAG9ylhW+HtLuUewVkHxlbOVdT6BKdJY2wMnUcZAJd
bCkyaQrye5xhTrWKtfCIdaWkNXZ0Cs2kb9HVMLoDJXZIhz3ONzhCiqw3DLkeDcrTBDO41YJ7xKFW
KWF+ZkCvhHsLpsSTMt31bcu4Q1K2Lt7RcK2xH8ycngLreqIeUcHdEF4djv4jZtOkhv49HN0b+qli
IhBOlxEqrtFZACOKvI1vT9t9cdbo0djhfsIY3y5ktCZn94pcnaYRuVRKWzE/SwwDhdxLDLNDEYPP
JkDLRJR2F6X3hThxuuiar9JkEjxIiUimmYw8ieaWq4mSQd3kJZLAIv3v2ceYnRmOq21qsB50/311
UYVq8mv99tncXF5j3WLf8WCgEoOR+GrJJhNFHDSN8n1DXF4REL1IPAAwRZOKnMsDOXTZYBSAhiph
Q0GA/ZB3EAJobVoNe8UL36r5ZcQtdpSiIGvGYxRLLFqOx/9RLb+hRzzMcHb8HaInvTooTW1vezja
Hd+M6SQP6Pk0hM2/hCOG4IoCQhrsjMomp0b2mBHojFyxVYgf/4Kn9wqP+KF19yFqfEuPiVNMmeBh
0bmnsyv6gBriOH1hDCm3B47tQv21hssbck8dfziSeDNBirkprvhaXbjnnHWB3baFhHndf7mJ3fXe
J5EM3UWQkz+WUgtsq+rQNRIuW3PukI/b2IXdfNXiuzVJBZ10b3Ya6X9aIOp19xRMgrWpqeYpotO0
J+ATE8zl0SY0t9eUTNpnRzrJinDmnYj0vfWD0IUjnyhu4c5dH2ntyrqsqUUrGJD5XN0pO5BUCazC
rIbg0Z6+OVhWb0ZL+TUe9zihlsrgUPn4pg7hNp22dGLfME4zG5YqF/BRt646fAeuh16JvSZYExKS
9wTUDHvT1QkQUD5n7cacuPN91CHhO0fFdxJ6TUyRHKPvCVDSlidLB0onJnsO4PSstivYil8XeQeW
GU9+b1DwA07OJg8Tli0ocTdQk6hfRyKfquYVk+jS8xtcZcs/P7uqBi+JcUWNHQrZw6MSSvvp7sda
0lwmYliJaASyCqy7O0TT7sHUciRdf+hbpk0YUzQkpa/fscHjtlLf9x7ipah59N4f7DqVyQlSYB4J
6ZC/lPn9DVZxFdRUkGgG34hutbNhx6XG6dTYlNJMfq+c07PQ35wSTwxVKYRl1Sv1zyIFtohZTnp6
20RU417qf14YL1rZxbhLwwadY2xY1Zxd0N26Msc0wDW5a8LIWOl7iJdSC0H1YdcWiA8vJG2TE94s
bUFG/BrUKaLmaWFDvd6dSHDepu9VLwTcfitimLiu+JYN5X2yfP18caZgfy6kh1mGHXSdhVFqvB+l
Aoyj87eWE4yH4dmU9b9ld6r3NDzcyLZ3A9LhHjL7ttPKLgzliLCnd9G+np+4yG7BCHkxq85n2TTF
TYDtwc9rJfHrsXIcdvW4XZ2a2N8GM+Riou+WLGEnUTM7D07Dt+wqEqHUXgeWIJimhkB0z9R4av3p
CW3aX+Ppr3mCNp7w/pi+gGSw3v86RZcPxRnchehvyED/pPog7/wP2MLWzmXhfBztW0L1DHah33TV
Vr+yrQjhHYbfaNEJesZR+GxTQ7jUi4zOWfwI3SBrU6jtHz4iHq3NlgTQQYFUYHamIgvPvMWFWuap
vL80UZJqV+m9w3RBn0GEbhbSSoZ6D6FoLZ6f+c2r8dIOfa6+4tm9NXFKimSiUY/YK/6iSJXRnK0S
e3KtcVYMWTqdDzMh0D5dZSp8hRmDov88gbnu7ziPZANHAFMn5ORPZoE81f+ypVLar2IvQUoETmVm
r6JrofqxIRuz76jJtd4Bne2S4uiHDT051JZ2BdGborXweslgM/mN/7v4aDcl4i3p5iY+CluaeahY
bQoilQ8WMStmlnFce/+c211gF4pXAVD3+BVVg6GspS222/J4cpRi6xX2PClwpIHcmJ1+bPAE1USw
mS65NkmqaK2dQ/hxhK9BMUKTrZuWLemC+Ofn6igjN6kKYz4EkUN2wOGUVayHATgVdi39xdaa7l5C
Jd3xe5jLuVlONIj0AcdvPz27NUFrBjAFKF2wj45tt07COOMVkecFbcX4ecUDPHSK7DVX+Gn7W5VH
CYwE8IMideabWZgZyuaaS8+3y93DXoJ1MY2u89fJ5h7zkRb7IpofDN5oTpH8wwDJi5mvhVmSyeJd
uTjZjgqjo3c3xgIfT+k8Rkq/qS9C4lzku2fTWnc2WtP0X/6eCT3pgeeHtWdDzc0j3o1V5wwaovd1
AGElrhSXZG10kzULATs9g2j9iw/e6iuTvPTh3XmUuU28HeofGE8PxlaWIfFpGZIyAlxGDLspB1ln
ymI4TwgwZ8PTy6Z2bQpYF31JM2VTWAAm8z6ISCujnqCgDLyX4h6hliOrEP609Do1y64Rt0qTDQoW
8kFynAEyCjaG+k3p4qbgAFwwvDw2lRMzRxT2JaOprC7IduRwGBHJhb9B1lwxsolssE5atoDuRE7s
56IA3vqikbcERIqVsOfZrmitnV5pOJyCtSat5hTu0t389FB8japhNjjjNCi3GzLKw6dou5x+C9D3
dtDElfLCnQ9XVMEad6VYBadAaJqZUo++ir1UDAPG9F0ATas0lCSEOwpEuYBGA7zOoAnRRc43bDvE
+2okN926WBU2qhUEVXwyW9Ttnq0AR0EM9b9/MQBoDRrLwNRRZQLcckPOvfNhd3uQEZcTAcaNTkgi
kWipJUc+ehr107/w7WXFLqlxGK0u6A2RB5QsLUzMfRfToADOa3X9Dxmcijcu0Rn8UY6+iFy5P/CO
/xN7cNtbQkdIEKl/yYES/P9qm7oFOW4HgaW4cjAqD6/zk7zEBGdxAxHEwGlUDsfYTbTmQkmWFDo/
bKmpZqx8Fcbpe39vgdeGz1WARPvTa/cxGGeAeZpAcUstnxeqmOQ459bSutcikO3qYqloZ4Cm1FkS
nFbpdVYu7VRLDGX206dvpkOvvoCvI9GYbWoSuieDK6IrlAl6+gwcNDU8hoz/eDL4j6H9Q0YwTBQF
h4isk1ZrziWE6zvAyGT22MfgP6LZz1lyCZsVHlweuqf550hbDriqiIc0zl3IzG2r21CXltEl/wt9
fEl7OJHTqhoJEriDLmyptX7885eQdJ/nULIUssuJEGnIGOzW08pZiL8PNgShWlHckRyOtPugakj1
3jTkXqSi4KpjPpquaDmpz9Wdqp1w31AKXDL7xQoeHHIkoKVd6JIB4lF5dzTgN9wf0xYjLQdpxCkD
wwzmDgZsLnWzmGGcwkmBGkm7rWZ2F6CB/5S4pzkRBbhzw3ciiUdhJFpgl57wIPG+PbhqgfErfuON
fjdNkI2Qd6H906zdbet+d0Dd6RbfYMt7d2R0XTyrwVmr8njWxkyUOv14ZTnLnSmjNuwUzeW+BZyh
PBpIXwq1WCyunkBxwb7eXfnvtRsBDFtZxSmV/7pbuOkdJCKmWHE9qfH0pspYNNdLn4dRk5qu78VE
KGz0ql3RhLSQqGLXxJba8BmfOMdvnZkfor5Che9wKP3DlGLGgG0f1JeeWPSc7X/e+Esp85tczXgB
CiO61+voXNNkzhiRJkks0rn2+drS/EAQHgyeQd3lGxAiGgaWOiyZv1MpvwiFge/oRUj41v5IRypP
i2XblYLcM6YAK9jnU8MCDN0Itx7VRIylp1XN7vAEsHp8X5zV1BJY0ote4kqNaWc42KPAJ9mOMffp
YwEjFe1I3mHsUJ0zuz0V7F3cbThvsSJdTGdXUUjqzTPVaQiXxhdDhWjVo8DxbomheAJV1DbHFN9E
zCbQzJ7Cpvu/mlp+iJtaE2wbgO69w1a+3cNlSUkIdqxRJP1eR3FOMc//qV1tQVOsvJyV1/GrRrQv
FYcuqQ0COUmgpRHOiDiKm/oBRwzWXjYi111sKTg7zQ1vVmIh0PoOLNIekEmVMAr8cFeBXhy4KseY
TUCxMeGBMfBUBnIH0Bfv3y8cGYz8C6X0GcSEkfTZahjqKwN+4TPOnF2IoX6fRxo/BYqtdnmZyag/
x7F56YsJjQc7tMXuc0e1ONCd0gwfu3kPu27SefEwustViTvRJdaMemSOiGVQEt+RAXKdBXj61R4w
wdShuUkZ5l7kxRREferKoxaukeUHtLkP8cl+TcTm11jHxPCQ+qfucvNUm2I/77Oph/QRtfqcg18w
oQtzreLsNV/LaYoY3/QPb8qzeFPWKCKq+oiAp14/lPWX+k6q/AHxbctKQ7iZTY1SioyGe82yb5lh
BQ26yqBQvbYv/xzLGe1qFiiyeeH+c03MxIsw3leOwBcDRJR2pzi6N6/tLFERAggFtRHhP+RjSRpo
sE7QHe0onBHr/rTMy7Bcoott/NqoKrU0Y8SXP/X3/0mZxHYzb7JhrsQeoPeLl2lXgw5mG9ASgSmI
cJU+IwvhEa9XnG8zqyC7aD+wdcotKArayTLgEnXYRHFCuNzN2FpLTKWCeeEZ+Y672hPYa4vKDNRs
bStrJoaM8HMXSNK5wKTEiO5E917XxBBJ5b4HCroVBbGqLZU6KAPLUTesXv16fymMyNMLXAHYfNC9
0b8ftrxqoO9rQ+bvRcF0vxHMPHEYVOKj4QzDPCY7PRQ+rKM3FYnxTDzU9pr8E9Xy6hmQgWzEbC94
uNQAc/mnI3rSui1KoV7IQLeqqTNp04QlckZizo14PweM1k9n2tiTkh8uChV6q1GZEotKtlU+qR7e
l7pXMd8KDrMOCgOSKF6cqhGucKxQ06zgIoapeKahOp6nlcw/hnujCqvCVOuaksXiX8xI6+v+mD8U
6bm+ik10yrhPFWOs+VmU6S0Twioo46ODFavSHQZLtF93A6hIMgUFqfmOB0D4glvp7xmRgjxkaDy9
oaelKmkinQ10DzwyzyI00+ToAZOYjleDTnawfOKIPw7MLkQq+c8M2jDnYtzGtQDRHxmjJer2eJwD
FGTAH2Pu5x5rxyIvVrnL9PXfZ8UGL6ztZE3jZli1EHlve4qHsWg3US1d135+VVdCtgWWzBdN7avc
B14HHQh2KYgKPYpxR7vdyz1VUiG4Xw9ZwV+aeSJm2pJE5Q195BRwOYJjd/PbR722/lYSlf4n0pU/
HmUMoKiJJqSYdSx0SCobbW6qIX6R4ec/jG9Tn/BVi37OZVEUc3yZV3vsTog3cipPyJ+sraBXByVO
KLHRY/wGbYixkAtkqvvBLfG5CTvk1FgQIp77Z1JXR6Od63BL6AcNNxd5tY5JZt9rtoeAm+a2jTco
3osRx2SPk4vDylJIcmeSfajgVjw8A/LJEoVTV6RxpvLblC8t+yZ0rVeJIZRa/eZEyCFXUD9tY/bI
561Hyz35QepCANrCd/LtCAEBTe9kZF8SJSUn97T+E8ImdSZL4xaVTRmP9CzEnBcSn2Ah1lpcoyAN
marmO40ZMPyOJGF2NPzoaQnREL7J0CZqjRc447OTrGkXBRz9HuFejFRkX9Mv8Fm8pgmUI2JLbYcR
e4chLjOsyGXdUP7PIl4TQVwaHl+0Au08GwPlq+8MckFbMiDI3G9s3a7ZHs0blwyVsp1g0Fwt9XQw
6bZpobDLkGB9ousriEtqqgLREeJl5eu2OdHN8uWXo2xlg8YyltMEuiNrmbrOZK8PKhHi3p95tZuh
23rqGN6MaEj/C6e0ubLNrN73B/RemXSytb0eBAIPhor5ncK+e6vRSY9nsiw6TQjH30owzq1RESJX
7YhN4W7hrcFuzhdrA5YEUtpOHeu5zJ51avgHKpgBZD6vEaRx+bumN/Wjq1f7SBA219q+EH/JOtwJ
OfoAoJMJp/5oLeplbgy3Ir4pjSUfSmBtWT2mXMsxk8hpV62GAcsK9SCZieGKXh/b2KzlOZ1pvqse
rzOZ7+zNBEZwTVhtsQaNb+Rhj6bonJrGDtUNAYRAQW+z9ov1J9BD+M9UGBxLbfxDybY7NV/lJE2z
iv9F3A7dIOlXjVk319F0L+z9ZzOBWW9gF6WYEHifmjyPu0g+2O7TOijYtiux7y6idccZ67Fe00Z+
unXawB6ZoBlmohsiV958cxZvQm73w8u2SMJLljpdqZNsGq+PQ//aD1kH6x8/37zqXaOEpU3tgom7
a8NzUbOqH3FbsDhXlW5DjHaaFuH5ilWqX7vWjF7wiYM/McJJamtymG9seefE2F7m30fbo5YqfIEM
GaD6g63Ug9/Tc6ZY7fgnltKEY9Zx2+O4f4Hs18gIGx95Omj8LodAD4tV5aHtTcY70cRyNOVBfc+t
JRkqqYfSwgdyT5g+4vjvi8wYySrKKe785HfHnFZN6jjHAr2OymqL0t2JjL1T0DH/UWiaOoE2uYye
oOChT0AhOHIzGcUIZjQqoaWs0Ftvj2dcpZT7wfz2TIo608ciLTifW4NQ3Q1Evtl9JTiVVyPgbApM
LBxu5wSECg7WxBgKQZk99ZiYetIf+TRzJtLicYgv7fgkBUxEpj3+eUv82y7qIyelRSJZuznCQFas
Cc3E2fm9QeGXUjNueS1lFyf8Y/nIx8T91Rqjnz+OPmICUIOwjOENihzgpfbc5Jd8xZW7cDaCeuGg
up8YXPqCBziwiIyZmMtfib6/ljCCN7cm53QnOPmEztz1JBniOBoM2hoRiaIgsbniejV+mk4yNTX3
uCfRjGiH763i9abXJD0c7TajIXYMLhT5FB7jhGmvsuhNfd8BazDSV5H3TKZ1OJUF6TjmQ9PEAN4N
JEwDEAG07eqzjXmWxbDm/XfqjfbpA63DNPYHEe/sd0mPFN31RYO7DSQD4iukROeFlRd03f2imbR1
p9xdIxgtad4/eL40EBHUoQmjtAkfus4BcfOq4uz7QCdih2agtqY1Tfzt4FlkTd25L7rkwSVWGgg3
cdSdV+9s1eOgKpXaf+nBgKufLA+RywfFH6IKCHVeGrdSRT1QmNPNg9ktS2gnEW/QIk/hLuVOK3Cx
1Nts08J3c8mHl0ZXRaq3ocoJIzC+EemIXz6c2NBpXXxGFYxiga53zasWVua7dtfTOiAjbgH10LQp
Zb0Z7FaJVas17mgiZkGWdcQJ88l8c8MRfW4uyl7r6H63ClUSG6AeoQSk1tJkjK3cuWSjnZCUcmy/
GMvEbOlCsUIsNT2vuezukuzPzcFcg4dcyOtcNUjOhQgoWandc8xwrhfSd/sefpq8uLL0w84QfUdK
oTFD9rtVQVAOx01jy3Xv6KQve6+RAx17++T2ebz9nx+LplCM+qXBzjPqhYAS7kXIPonsgUpjcips
vH+UXk/npBfDE8djixlnqPkjHWiyhK04rYdvCqyXrP5DTmE8GOjxu73+SXkcQEZdI5UzsktF1llJ
hwVVcwfCgcaUZUq9nEVCEsF3TkSvMoBawVTVFnB6/GB29lIVUq4KiBcUpNSQcIHqYjytXSPJe17q
aiJApCAM7sG/bh0U1CkS6sZvG64uzu+7lQq3RyZpKFmJdRgdLrnJBl2imv8jBMScSerzamwK8FP7
Mz4C9RbX0ugUcqEnEiXq/5uWAgMYJWgnOvWfjCM+hAczS+sQEBMoGXxn6UQ4/CLjgPn5+PZEBc9W
nH4NM/vE2xPYaG2xngU7UUu/eZu3V+6QuCf4+cPs5KpJl/w7cfHnZXVDbzD0hB7K5pwHlZo7sOjn
OhIxpeuAxbIMmvc/PVvUEzi9WRQOczkPJo2q99xGFsr/y5B7HMaNdnpgoQV7JAsXi0oj93EyOPhL
RxPS6o3RftMfhdLLUcomDYrwwhGAGP8H+zoPBDzbOFi8ubgS/ZJmEBV2G5WiSxCGmWyiQKKlqY3P
jMsyhqcynb8eFo7wNkisX9imvX4rLTNDaDUkAls8QyXCzkWfnlSK76xTaw6+cto/SzrutdFx0lr0
9VoNMt30NC/tHzIsp9OAd5j5BjSkumUQvkdxJdLbB8Y/XLKsVQPvpMumR0eD4Dm20gMvEB5gDApc
XaJ5T3uOi29uAuIO75a38rUhEJ9NNGHVcIduKb7884xWFnKFiC/du9Gz64VRiAM6534PJxZ9skjd
JDwpPmLLAEbypmWotyXBUr6PzBSsWlb/jNypzlTCWnTcFuv7CLCt/p4JXtPlQpzZ68/psMAFOEl/
gxw6Wvjcj8HPRltv6yccTG4zOa/buPXSdB639BAj8dyprMhja74+iTX6DQfEYzHauo/qDEMWQ9wW
a94iOE8yWu2EZJsPz0wPlUpKqR6Igl8RhSA+h1rq83w3qNaW9Uh/WGbxKs+xlMq7EbsVSxXBeDbs
+aNsfv132HLXnZBzEzz2lGoAHpmQsqN42wkNT4nj9HH40dPNuzVmJxAH0KlilEoWbnBdoUD5cAx3
2Jx2w0ZzeTvPWdf0znqBd9sOBCtyodrrgBBkMK7Rv4ay2Tf8c3KrMtNMceVL7h6umB/Gx7SCX6q7
k/4gC3QTMAC8grLkNLsR/WXctL07bKMU2G9l6YaihYEGHgP3PhKDna2Qw7/EZ3Rk3ZELEvqYGhvM
dqGQriv3NuUnkgEU7Mw8iI5u7n5+Sw0zq2ScY9IGff8LKF4VKgIm/YijWI6hg+Vht78K/9N4MV0r
uA6XmjEBi7juJ9RL+uvIeLumiCg+6t40UBxo+U5bMHI2K4NlCDSuTYRiEmSyav9U15xSfLpGIetm
XOH0d8dRonna2pHPFN+FFS1rrcHorTE93qjFKpPipU4ys51aARhQIyRPr18aDQ/9mkdlTETRui2Z
rWZ7JAVXImjxLk2nr5JIiQ/V65CdbGXedq3Z3YYD/DEfnvtuFck64xwDK1DV1btUSKyHgQVkG44l
UHeacmCJ+li93hvDXnRMx9ORGI+TIsiScilC38aEkvWeSCxHC+phTFfAFAE079x7zfIIoj5mbUUb
vzlxMdVKNur60cgUbyX0OTyn1MYgJwNtACbUU0PwvCFvxwK5e42d8UQUKEICrcW4enjdM5McCKmn
4CxONJ9+wWA+iKxKQpM0FXhJMyuLe8+CzECjn6jpgARUQRzs5VOxEJo8B6FgMvKk/M/bK5GjNRZ/
V3+b9vTMiMMkoTzuel3BoILjdmVZr8GjmK17yKb3StWJyClbH/gpB3WeqV8OFodFvGWAOADRzF5V
wFod5onOoPZv/mxXj85FirKS3YsQGGGCgV6XC8EVJQ0mYciN7sCqd2BZDKxTqqcvJBvtpl8t6U7n
pMaiVzaW+Zt6akuaxhdMRedzqvKLDAkN8/KPEslPAWsD7RFGt7N0v0vYcX+IVKpBLi2KOq/PrG2J
oWGpvojeXrnYBd0eChlIIWOqZMMRMIrZOrFYliLdeVrUpDUwN74166sqyRo5edF6+f/n6P8jANJ0
qlBQoDBQOAljb6D9xRuXrZLxQZHM7xoAOqpUgK3cEYFESUecUbHjx4V0HLX8kjLBYp4fyUdxS/lv
Y43A0dhd1yQWajCd0YsGitNj8vLvdISG+sHYyFcIvgYZhoIRpFDJSF8hDC3+3fg1qrRE147f1IOp
KBn5KB3rWz2Khh5ou7wWWN0y2rCtEIiKNmxAKFMU7cih07+tUx2n1tGMJ5UC+UGdMB+zjScG6q5I
Z57sCAvkeYA9ZjXho539PLMv5YRAKk11iXhZ1h9ODyEyx1mpfujaLMLR7QYkkww6Bk7n8OPEU3wX
wDnnAqUTh9xBDlBJW1bvrQ2PTxbgzjA2kpTNrh9QB2t/mVssOiNVGP80NvgN2Ekt6Q1a2MKR/8DU
htBji7ley5CQ9HM64F+QmGfHjpZVCQLmdALhnyqIZvawr7XwSOBUbOg2OSRxuIcmAxKQBlC0tQR3
VEEcoxmh14C/xJLT63x8oIg/SLwtCKUXs3vsD9r8aPGnUMCZEVaVd8q4c7QdZE8yeuwqoJYEGgBR
v6c1QRJhFMnPEc6VMLZhVcYdpG3YoilgFJkaaLG0anRMVHiRjumbOHgeFtN3tNSSxpQV1B+V6nyk
TUEgq7f/688lp6itPQoUbZ2uSDdLUo7Bt5DtiszZFMNRQtU3sM0Sb6vEIKHurgYbNjpzV8EgCxw5
v8mBinC5Riy8O994FoASgSvx5PBKY3PCvbnT2o/26rsv447BvhLUMjRyqRt3WIoKrDw2pvIbDGm3
THLYqzsi9AvPObcyvh6/fLaOFG9fncYWZmOIirzJL3yb8dTkBptlfq7XtaS9tILUuJRycmgIrmsL
/4J73tfFxN0i/0AigAPGiYtpcRO4T7Niy7u8RZJ3+4YaRRWcJDpAli2dhlQogZYZPDchKUibhqTt
se6nsmJTfMzLJtLHGaIGVZEJK2Ba7XmxUjkrmTLT3ifDbbCreFMMfkYbEWT4u0BR0dKqjyR0JWUz
zK6yEedgxrVtS9fe/rLXbi0J006uQUIiACkAu4kqyny8rdYdeOsZGTO/6hBTpx90GvEuKMplYRut
2MG0CC62m67VHNFwE4IYDL5R7nsvkZQZPu6q+ihzoODsGC8L39J7luTRZygPvbmZ/WYMHdpNbmkp
KKDVYZ17A5PkapFRSP57ZrRMEbwyvdBzvD7YCD4DPBJKr8n4R07b7KnpK6N06bF/OsrJu74wGwFr
uph8XiqMNgGqPdXLoTRvu+WH7LXOU9O29s8K0DfmCRlvGzcKwQCralUbMq2MBUScmkRNSve3ZJ1m
HheBRVjynOWqQT5BpqAfd4Gs7Q9jVDBJ2D2AbdSxiWM9+rNM/2h5sNyMkx/+V7u94NDaR7qhTsBO
lN6s2lkm8r0qN3ndwwfpG082f9JZTPEAlAN41m9EQOBEDw+F8PWlXjJSF7OE/Xb/63gbo2c+HmXa
4NPCA/EDYXr3bf8mETYaKyveX/NqUwFb1i9kGlkypXp+0Woin41bFZ3EDK9kx0x58QaZEKlBUCFJ
XcFDMtLMKnebdh/ZEIySZu74fc+vLx7xsm0MRBXUnwNPGjcljZ6FCjmpDf65jloT3Svlz3hyXpka
Lt0By9ZGWzcVRYYDUnYF5V3gXl5L0eu3Eo8vGZLNcWEYuu4CCe3RsnjqLlsKJbL1mU7CH/5BUucZ
gACR19EgddntD3/NCxB+7qUesSLefJFFs6yHYyM5OBNdFhJ72SN+wKLTxHi1EI4DNk2NNvv7P7wg
ZPo3ZXFT4+t8a79LhBnHy4xvZcZBQsYYHiWnqVePZhesvT62eS04qr6TZuvwykfCcSxSM//tFZ7P
odEr/oWM/JSdsMYLPH2DxP49dwr0VWDua/kqstqBh0ryUmuqtRVX8Vwcp2VvVSiX9kRxjp8lqCnf
lyvqpQ9ciXFYZbtPnQ3jZgsfKarscZYluJ5QsJr8ew4QWNoDB7I4fiedbRzrgYi11dTFVds+G58l
f7qo/zAXx2Y/AUr7BGYF2RP71n+b5b/3D5ry6Az1rPO4xZ0v9qkMYdp1ut3RY0xUEvFUTvhwFcnq
vidAsawS5gXorXJ3j8G0dMnvPU88twsmE2ur29lOU1JHlddx6lciMm5qzf3uIf8b2OsYXqUC8btR
hiGJCJ6JEZk3/DWoU9OPbwRzLBZ9qi68R3XzYOZEhG2LaClfIcexGN2fbVwySSRPtAjpoVr28cZW
sdabaDCMp+70JY5IlBN30w9B/NXi2Fqd9E7O23h2i9dkXUm3tAyApMZo5CSQVPH+aHZlTKjHc6O+
6us9LdNHOnzVKvtRVeQuOVDMoLfAOc3xMU1uynNtsTHrlR9VwqFw2NbA9jR+/zx0CXSagBu3wVhm
B4n7jkuTtUY7EFyjRujzwe+YwWBOxJbm0sBtJziDT69vP/ULk5Y/t9C3YhpCXL7XdVK1NwMTCfb3
NU51P8bHcLQBEjucEVcWCmP03LqIj7UR5wvSYjBRdBSoVQKp2gYI8s66Vf0YXOZVH2vxjFMy2CcC
Koy+ozC7lpBR62AcJgv08Rt+c3wayF6i8m8wCffVhSCguCw3qUYWU6s7yZctHOoHpJ0/xefIy6Ca
FNRVqHIv/kh92Hc/CB550jN029cjHca1iaztMiOl3ZsZdVYensFkqJSHzx+5cgMSdF+lyfTLzhUe
W6hmrhVv/5v5BqAi4XfpgNJnYFjNL4PYbbmBHd6M17tyZCg0sgy7QpwZcj1I9Dyj7JxOHZVTaC6j
5smF3d6neoiNStrgYliQU4e+FobfN5CVfJ8vZYsLTVtW9ZBCUWdj9Z5L5f9kJ4INiy0LfRGB2y1f
nuN5mSeqZGNNw9SRCC6XOO8DxztkfwPHUPWAqD7WxN319MOWYLRmQab9SQUPP6aUwUA19/mwRfpR
ftyGsB0XseQs4u1stC66M0a2yMmdxfwhc/H6Rui98AjiD6qD+WULg39hSAO83Pe8nvD7/n0p2xnZ
38Gxd1rEEMMteS3RyjeyrOGrR5fDY7F/bVBArRzYvBuC6CfjCIRAVnE0AlbThV6aS8IuD4f50xlu
aO1RF3UJjDJdpSjGxEGDm+yRMH0XNBHgPIc7Skmk26GkVgC5BF2f8AmutyEP4DKENevOeXNq/hyT
2Iii4x/tnNB8VayGH/pu45quFOcOcRL4XDMeU+D21iOcSi379+Pfr4hQHGICY0Gb/55I6jh35kfo
0RX7CQKgF+NQIJczltBc9VmGeKo3K3QKHy1b3F6Jlza4rCXjhhXVyMI0jpon37oSlIiQxI8GP77G
EFTBQWLJw3hfqJE7GVNeHS91et/KqylGvm1giwMkhbSjeLEw0O6ukF2hGB+kVMzcxmHSXT3TZzDr
a9Pow9qWVs2IIqpma/ChuRCPaZOUbBygadI0nGTLVe2L768nCc7w6IjEAl2/qZRQe6CuaEFZlw/L
s3UO1BBD99p5tqO+mB+A/JKE7SNqNKJ3+Df8Mds40Lk5Y8M9nTz1IdkM/n8SWGKA9KrwLMS+EjRn
RL0MThKC7EQiJ5sRaQDueDu7qCECUjepCkIjwyOSBnvtOSo3kVO31VeB/7Mdvp6l84QrBnX1oA39
Wj/K9oY/v9aOFjcQqGgGh8wbMxEc+vWbLj3RRH+4JXtZtMy2oWyxFr33Mbcg1gPs/V9HOgL9ZB5A
ztPNbJs+azOBbnlNK4KsMd7MPZSNtGUReNUXeFCmQfwkE4dQ75YEAf+sXwQ8jHURLSK7ZEVAVg+v
PX1zsllHK+G3APZArjfuroHyXSKY7k4lHvEjp5R0k32hQqPDCbx5KyjmVp1n4rntis2593lMo/gl
OrUnIEJaGyGdophcC8jQPFDaOkjLakth7cZoEN9vWOXCVKfmFSt3n7txGg+g9JKpwmHdgAI1bidX
U/fvS0VDUPXHDtbUzEcgoY1wHCibAxwMz+dIb32VI4bkBy0205/90DWPTXI7wdO8MqwlfFwxpJiC
7VW5asw+YiHd7dZQaRwAkhKBqe59RKPG0UpxaAOsmM+QMwrZJ0x6322X4OjyTXZSc+b7WQu8vKhG
j6OI4h6EnjdcuZmhFhb/204hzbhStPsW/MEtwPKEkC3E6/02+ASdjl9w0luOgC8fSUKtSmd/gSa0
0eWsuV5YFGOrAcxfEo1tOdOH6xZounCzGVO0LSpJsrwKfpxXJdZzJ8vTFF6aZeL6Nxmbc6fQnbRF
J/4Z2kOJkyIRVHK7dDJmO1SYxzevUyEZifnjY9C91iG3I9D/0PWH8PC2Xa3P6xdF+7KEpTha5+/5
qOwEiKNxZvXsHfcLebsHdlGfAHrTHrXWVwjn9Qe43u4/xhR4iQ4lnlB7i7Yvj5XG0Tbr1KvHlpUl
6+/G2tVqUdrFlyhnqPn1V8vOM8uymt5CuEBfW5MEyjPZ9mqXmnQ5Sjo6XWrSHx6dFmHa9iQJqN00
Sib7Ppdot1USZlvPh1vYSpxwB7epv8yQ00NjVbQwu8EhEFf7F1oo5WaJ+kUajgWNeDwFZTftbHi0
MkWv/sBcqXwzQln2Cxm09TWSUk8PzVmNXsSu5oecJkqkXz7g0zJIGsnDKbw0u8uVtjinIhNBfFI3
UDsy2wYQ43rlwPDiCkhCtAE35Nrjp/t265t35D0R8CZqDYlFO+XbaL4eYmPSwO1HiI+yqiAGoUru
cLvKOkUfKuxR/NOLks1SHGQyxSEceedBcq3NkrIJUCiX8XJfL+Cxowpi8tKFJrRmFRkXYlhtniN2
r7ElaBF7JRMctXbS4kL4argpSjb5Am4eycw/DiC8HaFnOWPKLNqU/8T2zzGxUHaaUNvNAR2u1MTb
7KNgsQYk8gqrPCyKehv14D/jN8rzn0m6JJTjbXh822/yGBewqZzLpNrKN/IZoV9OOn68cM9AwYtv
QqMFe+ZVDp2hjqY/QH3mr0iWsk1J/SqUmooyI4K5j11z9M4Dv07THf5aqq1jFjJzeCwaUmGYICpH
RpDs2EyVmSZP9Brk3nKBoGey4VN+ONJCIAl2G9vmUS+H5QvRe6kpuaW966pWlr4FuEcQGa0UC2tG
AiO+Qgli2mXzei7YkQTxibqyIGTf9qA/rEHksjQDP4poj50JvBWqaWMETCzKwbOo0aKh/5ELnX3V
2SssJnUz52pWr535JETtbzp0DcAccU8CuPnQFBUzh/ht8L/2rhbPU++AUmEpuf5uEuP9By6vPLLQ
qXiW2+oN6UuPUdZG1rHHYRP3HqMw8WCOTC8CIVqQKFb/99VKUczWtaUG1wZRaez5FuK7TVOBXm4f
guzGZK6vdR2t/ZOwysT01F7REpe8eAaNKSUikxb9z32r9Dy890vQFLl3+gg3si0M0vaKO7f5U4j+
C+CC9myk6S/xUjfa2BLveKiD5z3l6slrGFZhHSmMKsr4FpmizuZdbw+QTDo9zRhoBlS6O0FAqbJJ
D6kin/T9x9HnvRTZyoWaRbhDV5c57AOsE8Q4c9AWXLQgLVGfiwwNsFos+rqsR+AgSn0TFr3n5fYL
zOREsP+c40Z2/QA+owB+T1ppa4PCxKCl2t7FEZFzxTqKeVEatewykShPD7CylPhkT+JAvu0V7KPF
d8DUK2nFI+SneeXn8waJEvBQylc6qr6p6/p58josbOEXVapjgGm7kvX4hIzFy+/EccCLr8+g5cFP
Z+y9dalVYvSJ5fHw1GlmUuMi1LDIvReHDaVdd68I1a8s0tXuwg4XgEAseF+I4SlxfRYBtW7lYTP2
Kc5tTCAyg4vv3mnTa4o/xjq0E2IkN6p3qcGex2m4TBbO/uxSr4nfEdAAZEM5u/ejm51mGpxyrbdW
GS8D+4F2S6IY4k9W3rq2/kGogrgEzQqu/XFfC331YJ9LTUHX94XlUtwO72ZrDxIvRZkeKaHqcrUN
YPfG2XdNltKcK3YpuAhSlSuibmm0cXFy+3Omg23NoECDGXwxLyx8vVp1p4ITEw+k/RAGto5dyCLz
XP1cBuGc81bzadGzSAo4c4e0MWrdoCX1kaiBuEmrJBaLpdrOeLeDqIC+osktORwOMpIzweX0tSeI
lYjNjhzAa89OutKflQJ7MjidZWnMZtOpuxNe3dkIEy5EyBeS/GBNx6Gs1+n8DTk+LpT52mArpsDP
kBG+zLXQK4zqJD4LFiyaJk0edQ7FpH68/Q04RIAdhUw4xc6l2H5MyCbTEzsOzee7H3bNE+zN3DGO
C+ZZvRxHUVbPJKcKo8jiKvTToXYpX1Qh69RdKo8HMJb6/r33+XB6VZ5OGDvZ+3c/OrfeXu5rPJ/Y
B5HacoYXzfzsBWL6VqedFWxYA5qT81LEjE3JlL0o9Agqui6RH3gm5zODtxUDngcpc/KOauRi1haz
tvE4KhpKD01pnjnqsEG9CZymaN/ZzQ8yo+0jM1gtMGN4bNBIekrFV/AEkpEk07IqdwC/DcQueZvV
CR4wqKkcSP7ku4XOddeR7ULvAEqppsaG6jCzCePo74n1x2G7vwyPpuag448W8q/tiKfBSQI0DzFO
7HdEg0MYCpUePP6Cw1wYrBdiN+oIyYuGtWc5D0Gp9+ls4IE1ekLv8osk7XRTm9tTG1gQixpOx9JO
Lj1vYB+wJvEj0wM9QDpTZKKU1TjnLO22WrleuIIIoa6u4M95YpzJlq+pcUrm294FTUvZIl4Inqlp
A+zI+4NtEklVIiHHwGPpXfhtoXgLn1pdoZ1WK+WthqjP+Mm7W9XgCV4Rocgp/UYS1a2TrVwn1pVJ
dE8SH0eApUy2MzIF5wV8aF9KvbMT8/hBBH+T8s0S7Kd9XMrA84zkfb/etSjx38RMbrGFfX/aQ9BB
gJ2L4bktNtVJDyUuEI8irXo+dcDZ6ARw7k5NhCDDIb162yCFhL+7Ve0waoSERRZjOfw4CUvvxChN
jj4AOA8SY+0jmPf3y/J8GyE73oJEuVO+Q4mcL3sDx72XQYwjtUXJL8bb0PTn4BIkJtC/rSn5IBZ7
3HxIciCJqYpabcjVNENB/pHwkCh97d7qy4Pd48Tj1c2AjXM7aDbs/7ronG0sSE5Y2hg4NRC8mqU5
GvDg8P+pLK8xs2Lz5gllgoLFv6eC0YSbiYqO72e9Mb1AKnMbhKQxRS4GPs0wYjiTmstIF1IoDuwE
ue662k13jXdcPcRBtfiN1NzCR4NRcscNXqN22ef8ef4Lhlty6RvJmC4d1Iz9k64OQ0Sdp67HYRM2
R8fFXsoV6ewd3LuSIQj5s9vaRXTDeChIEFMzPtlxho+1O5BfcEWs4Xrb9sTBqTGz6V/4Fw6n3ozj
iBTM6CqDWylNoFtZ06ZiaNEMkZstw8f277uOLq+f7W+5WOLOnU84nEsGAhzuWnDOR/JnR6+/QE5d
8RAAEm4BdRidUW3zvQaCpCx2dJSE655nbraLAFzFS7jtanhfxawjqpxIhsr0gz16UyLJwb9tNejC
xLvYIQad36UTeEUxtA4pMHbsh7PXiPp+fG7mZmE2yJ9r7LJvI6IzcqCu85yfJ1N7LCjJV6DZ0joX
d1MviR9JqOjnFix6RuOLWUSWIPnRf8CGmJDLaSVVweb9ojciM4vIRs2sRJYK1Ha6nsm3GVkVQinz
2JXUwlrOuaRpo/8BRU73PYAUC5UXcL0YsAZunBjOshv1M+a1pM1gik/apAa9JoN3jdOSfTeleIyw
TZMCiXibejPy8SKJ6wX5Lu96tjEwM2+ueTIEjVEvpraBZqtwNoo8E551O9SnNQKaCDA7LksUBG8Z
2I3ddPundaAS6TvzCCC1f0NJfFSZKo9V3D8XBxJcr3YuQOSlYeToErvEGWZEV9RHl3K++ZUNBTzK
CtpCKivZ2IGQ+EblC+4M+6NvTxanPouOw+rwuywr/+/yVHRhZK1Gt+UO56KropoQ44txgzTOaHQV
7osmN3EdxyMI3J5xMl6NxDQEQEdHB0OFKkwJFpH/LiT/giWF4JEc8OnvFT+GApkJucmfbtIfzYxc
hzi+vMkLoh4msszSGItnmGLDAVnBOdvm+jD8Ow2G2A32eQ+hntfZuXtudJmyzyvsx+Y4+QovE1mx
l5SxJZL7npNhyXS+E4EZASBsRkeg5bRI+07i+3jCmufjiYCn9uS4k8RW+gGyvJuxtAzjRuT19WFj
xDQ6R6pqkenPCRGwnHmvQ3mIQz3C3ajrDvjzKH7OMzZYnqvC10PtTSdjHncGafnSITfp8YFsHU36
K9o5SK5y0arDNKb9oySe4W5RCOS3WOLQC622VXa30x4jVQvqe7SMXjmJFF3rTslIePaFVlN3ocTX
NxHuuCH/AzjvtYjgrYvAWfqX3jI8Eb3mJfo/tQqGEAXrMiiD5iBAgVsBHqUY+wkzp1Lj231YijDE
ZcV4cqABu0lM2U6YtaKhMj8M5BcdPDiVZl/Syqg5AOQv87+aMG93DzCy/QZCa/Z6BOY90SCa1vvu
e2imwLmOEzxmtSihjUAJhHFstK9HyaLS76zSUIqPYF9ZK0hUfLY4RWLiFh9JwRFROFOQFKfk/K15
lBi1MwYky/9LiEFIe2DeJaJrW+WsJHdKkBWxyG3xGwrWNKjaTKasHW+RmrDOb4w25U9JSEUOG+kd
qcruDG9RRWwgFpdsVvqPxFWr0QYfz6ZxsZB3ETdAzOPcc6UNLbzSu7hNwSCh0/OoMTAkzqjGlim9
yDGobn9+P41zBMLXIrKPHrJcLFQnSvWc0HepuORtgip2GgXY30CTKKxmLENIo3uje9nPnY0ipZrT
pAbyTLZ6m4F50gDhvuVqAHDeGG8N+j8TIL0MS16IvuSIcebs13t6NGKJ4EwPlMnNrJvbVTcKV7Jm
+SvSVd/eqvDVYjaqbEymKeIAaDR5Gx1dcK+RW7CQevxZN++cijIfADHfh9L3DZBw87zGnPxxRTYL
yrPbfyezw7k3q+atStKYVKREU72IsnqjoFjcH/3MMEjxshi+QfOGymO7u3tRusBcHTkhhj35CAjB
O4wQ7AxZHhWeqVJ+ygFpWWpcjf4ONeiJE7+HKXUnCNWYqL0mPX85mvNxaPnAJxDbH8pTVm2e2fB3
zGRnl0SOinudyLZXzOh0COT+sSj3bM1Wom8g9S5Bw2Pr/At2WzoyiHQqD0U0RKjojD4hC396ODii
g2wuW9tUitipaYg67GP/qYaPHLKiVzQmk+CS2sahyD98yk04tQk++gnjsqqgC8Tw4GAifskQSGvo
XyDcFimUbwSeMJK+QjbzotLei+aG/he9p1OoK7Lq29bzossDjWQDYonX/z9GWNjP7AGmiYEr3khT
gnM2OpQnx26x+NbgLxqI1lwlXZj1CEUvtMLc3UiBrWzKAbgAD9wz1vrgFs6hesJSrmLh1kjxCgEO
XYjAWGAoBoB556fVczeZHnZHcbsWvFTnZkpe6fEPfAgpp/rR70lK8dSy7sE777mo9zvby91K5NHu
4n8DRmJezis/zmNqJbs5UEy7pImSRo2SQgEqXroRF8vol+KxXkukOZyfnbKwp8nobRcH/juHc2Jw
hfmYOlXfmVusA/jaRRMc7V93EVdi+3dhLG7FZiu0+rT0HDO2K6fg+4p3HZbBgGYl5nrmp2lgiOvn
A6We0oEV/sqo68K1r+7N0pPfJAFclLqARC19IaztuUKCZ+TziGdIND2raZgR82s41YfXZDmUQKcT
aqT9q4feTZsE7NkjVim9zZR7GcLbYH5bIHAcWP504L9jiezyXYbspFGsv7rvBuldoPcqK9N9L5Eu
P+Z1nHlc3bTgh1YoTmUDeu0O5BghJfLKwjKP6vp2RrTqH3PLf3ABKMx60pu58pLMUoFEq7xA7fJH
2LYOnYsACW4+cqzcMjDh3LNO3jctdsfsnBsAd7SJqJ7QFvdXUYTyb/LrLc/PleQo7mGZBwjQYz5/
h/j2+tCsKLf/qnA7DDyMdG+0jeoS5C4pxLIAr7Us6S715XT+JIttKHYR8MuJi8RASnPVRSzrZarR
eY8q9t/kpvzFkWSxyC+pQRXr1q5+Kr7LcqHCU3p4kjiGAkkzgtl0pG34E4Zm7vyF6qecHI28mxdr
RJr1+wb3V4ywiXQaXx5dp1vnqODSDs84ndbO9EO551liQgxnI0+vqgMUeTEgKumPX2/KpW476sfJ
zDY8uazcfHHFiihkcepz7McXBqaMLg6tPBtE1xyC2MKgWJV5fHgU0UUKHSSAZBtPfMdxwsSDXg2S
rgY0H39o74etJkw57Bpz8qRRt9Zqz1RuznQy5cvnjRZFVRynfduaN8ss/BcsTgvtGCy9IMVfPiMO
QUKbXFQCdQHadxbZ7QLWKH/GpngpAY3c8ZqcJJciKvhAN4XSrZKlNAzbrexG7MQO3w0epC5+7VYi
keKbPodt3ELoTSEREBmGgKOzNBRRKmOyqsbqJERPWbm+bBv9cGQNe4VvkG6khqNskg+7Tv/QLWbJ
oEloGJnGFoNoMZpxPxECjnuDsxVYsCQJbE91/CgVez7vfCv1HnXWZp42nMTlqmZm/A2vbBJ0dKol
AqkOuZgoKK/mw2Nb8X2nPWtMTVnwIqlpI/NIhEumY3itlJcrl2BzInGkFb1yzc+B4SeIRen40gxh
qFaUcHDnssJ/UENE4GKQk3d/QpeIE5kBVKhnw/mkI95puSaTTSw8n4iG1cXEQJEAW/S/Vaii7UrI
iJQQ3xXLIhEakyPWZ+HXuwUUKW9J6n7EFvAxENQibQHq2M4fHA/fp4bm/MzfxMb02j1lvI8jEcp9
drKAg8XaTTeR002rIN5nKCOARS4xK4WuO7GUkAYMtDaeayMC6lqga1dXiklZgoJ3e8tPRAMpx54p
FjoEVdqQjhnQKrziDx1PuRnuOf2m/Sr3oNuS7PMTxeYhSJrsnthONIGCDcid8RYb6qnvny2K0Txc
zFqVfn7BZN6Wj4Ii6hMnSmTfmxW6l9UWcQBRz/nj2vLCyM6W/UIMTxWQZvNq+/XlorjppAPP81/x
glofFrJZtMsB34QZm0ymn+PM24X57js/lQYTKuRBS6KVJ7Mrj56rSeV0khZv0v2X1p+2E5Zqfnbx
O/NO7XUiCyyqyerxdaHHwV6/NmxYELY66O0L2RKWGQCnhLDk/4Ho5avD2JdjoFtFEjoip9lzukg5
LgAr7lHBGULkyCeOBfR2RC2hVawqV5zAGhyI+5REh3B2isgvJS7/hUrIhbLNC1igXd/W5K9mL2g7
Uc6lomaUv4Ak0FCc6f4aH71Rv+Jm1l3Q9dgTJWtmGZUeUqqastZtbrQ5B1Ckx0wKzS1jXoB7bcdV
66S9dF/7qTu+l8Q19TtrvYAuN0CEUiIY67kTw5B4AXINcva5FBRJbxb+pM09RZMVu6rHj50ZXZ3M
c9TMXgSbLH/y1S5Iunq4nL2rEu9psr/HCJQ4i4UvV5c6I6bLPsbgZgDp6k/+fvB0IKUOCErI6833
MU0jNLQnXFGc+Lf49KIkWYOLw3bI0RlkO2MN0RaS9CZ3hW8FxWkfS1vNAvqc9l50AaKkAR8toxbg
G3cDXZmuXUpNswNuOmnHCfe5S2MHZCjtOQDekCqJ+6dOE+Fs7clrb465QqM2hP+QL7wDSuube/4W
h18/Qf3l6b80+2Ces7WYP+sy7laCaq2z9wrEjL7X++wC6XlMY4JRLrTuG3mw/comRO05dD3i2Wj4
QuH7eeyAiCUZIcxyvETkAtnxQb+yTD8U3U6XMAo34cGcGCmFQdlcLYFMlmAy6h6OhpYfXgqmZMlp
uo9A6rby/muvhSUUIBt3kK5DKOiH4pAiPg2M2b3yFmCwJ2pxxjavx7rOcEGhdCt+sxhb/t3eZap3
ESM3xdor4CYA4raSdk4upkkLmTEmpc+Ug/bdlr6FabKCt8aeVPIfAwpAh1lNJs4MZWynEUcRZxkr
cogWs1qsnT2I+DTZy/aKGQTLO2iplGHxxdE03Xf/cnKlwtoKOUnJV4wEikdM6LN+TjZxhZnri52E
E0zb1g+eP2e5aq6bNTjQwIjmJBPor6puvLnK6rQtoVEMk2Ue5MRFQOZ1CkqAla6q0vYKXa5Aeyzp
KvdaWn39RYkyzba6hmKScTiHtmjuUkE5cSaz9txH+0RmtncwYsgKq+q5Wt5hlSoraSksngCr0BfP
Egie3WZ4wrgb1DUZNYIfKdfvymUw2WN32hBQ4DMXbx5C9i43Nn7mIciIA9E8x5BHRI8io9BqTIrD
xxV04CLQ/5ZOCpl5uaDKAMK1IFamk3127E7PaeIhJAP9hrg7+q2g4G8sFtUsw6JjJUis4toii2sh
1Oka6SWJDCg8p9zt5GJDwbU7Sh0xdoQV1ibehKQdAkkX+bnRweADgBxXfWv9xm3NATZw7FOQnHf1
hqO0xaApg7x923vKoIf0iCTtOKScPCgNBDoiuCo+2/DYojakcs9utIexJrttun6YmopRepCfLSlL
inQObx/wchQ79tu23fLmS/0HPNQJ801rbeMFQOZnBFcY/+aWd/BY571q58KCjbf0s0mCUMNdxJEq
15vhCj+7NuI+NNMJtaNpgxiBOfKeKjAFz5nim5z8GfIvLxv9MXubYY6Ba7alebB+UmzpFW8xjldf
ehM3t92nKBS11YYdyPAceE9fk10kw6bw0pZPaQfZhjRVlmaWZCuwDdGefzh0M5PqQeP1yVveK/D6
3AUtuoElxS7drWyG18sEJtnFSxg34q7HBAqw/i8xyJPzHLsakxVuncJDq3y4CWPaoKuwwEQjN3MX
MmmsJPQtdyqJ32Encqzj/+uNK2JQbymbxEAhaaEZw9fHgsovJ9zU+25YQ3XJvt8lqSlB5YOV+zQp
kXAMsdADM3jYBV9k9tDzRpjwre7kBROtUYIYtga2mr1JpSc5YTJQobR0y5FQhSpaNmoHGjsI+NNT
XYagMLbML7cek3B89Sddg5DTFC+5kHpAzzg+MIaiF+U4UX73thcsh7g7fV52HaWh4+WEyxc2FkZi
xyM+CBR9h1c0nSkbhp1Ye+0jGA8kFPz0m2q9aop62D7wWHKVxdKKjnWSteD6AxpexfPsa4LSRBfB
r7PrBhcqv+DPLxNyW61NTolKOmGjAinIv5p0ZOdmmMFq/w6B3u7bI5j4/oycryKZvmOYThnSxK1B
H8XdCCEDXkkNMON2tuvCWFxk4UH+CrF77OdpqQ5nM7WPFYuzN1VBDIZ27yKz6PxzMNPnhgUHe1TK
hc9UvVKhGA2EAAsuKuz7Xd8A700YPqFL53TKwBOp8qmi154HojtTH38EgNRDSoOcrM6Aq5eCVnCy
UACVzBeo4EksnpxZfvdcWjax8PetiqAZa+2YNzYJ5C4P7KTNcbPl3yrMwmJspCJtS8csAvKngybi
yAJfusGeHSZCZ4lJKXNaF+XKZ8SQ5XYnGviVB6uZCRPHuPadQMMLor2FVKg8CBk81LwRKcChUznZ
fQlxWa2N5kHP9lWqkjP2o1PNM0yWh0ijPrVZlaqMbql1tKAayNtrEXD1KMhVwriDg62nF599iH51
3C/MoF8qjC1NzwhZulIUXZY7k+Wc1Zh4K6T6I9eg2Nkvh7fdpNNI9QSbH6SYe5/5IOR+kQZQKKqm
th6Zijehy3ZUW3Hq8HzrXRb+Kl+aYLxV+/86jjgkT5+Dp8uBePHTzzUXgK1brjr1i8WxTUDK4RQK
MYfWBO3NK7ETrtcBYCJG8Q0J8e+JDv1iX1yuqR8FYQzp4yMS9Myf823ItVwqbRpc73sm9Qq7Mcmx
StPZjqJihUZoo5WxLKkWr3UB0udQHsg+naF/Pg0yk9Z26rQ6+nU3mqipN8NFT70mFyJRWKGaK1Iw
uVeFOFQD5Auc2OKT/e3ABlUYmI83mBOo29L8P82c5OL/MdN35RObd9HKkdbrHfy3fpD8WxFT02GB
+2SvDhiHYG36lmPqHGCRQ++T27/sH0fnUfHNWHNsc3IVbUrv8HuSMZnt9/ZQPot6HVQLR7NhK8ZK
NzICyKgTK0r3WjEKkL8wScrjkxC/LQ0dODIxwgY+pQdDIk5q/z4v/qDk1kQ51P8O5GQuxLdAQqVP
A+a7GMxULKht6hdXmUwmV7y1+gfuy8fQ99qXzI3kGdifyRFfXJzl9n9+DiQh6vcnlTbgQk45aPvx
zLrPU04xVPhwNllwdc/MFoZLzF97j1UhHW6BiDLfSR8XqkIoudzaLwwmGeoAgFWtDcIFQkgKJU1h
hKSa/Qa54nEvd8640P+thZffA/UR4lVoZMmZLpNpmLl6tM/G2TNGMf43NKYV4aoyfW/jIQhLrnwF
KbecrmVlg+OjqLxDzNlFEdvD89/NtzFmThQtmVRZVBdHoAXKJfvzbRogHWXXjA3RL2s1i1YjJqsY
HoAg8MRO/Wv7dkrkp6JMDZ2pFQ7NwKNg6RFJgQxY5jCTw8k4l/QksbfqyzuUmxfE/N1bRoA21hkh
J3zufQo4uyTTtn1ppAQvLnNggsKjgSkE2a0NxkAHejGej1V6+XG6nDzjUvWtyt7MSGt6D+KACpxp
kqaZD7Pb5U/s5bFJC1horq4j0gMvRAOanTwaA13SoF67eKeLTdThwtiXDLtVHzfT1X9gwLCuusQP
Kl8Hph+tIquMmmNVEqIZY85EdgpxLA+cfkbCIddvNqBCvDgUov1AkTromzZP6WB4XlJSNa/0oo0X
mliNzGT9XfEC9n4GP+mv0Z3P7PjKkz2cDpDAVilU6onHl9p49KoCRZPHlTl53yD9TYPJTGqcQz5o
PCBqafYK+dpBIGcHDqtCka5D3hMJxOugYLi070qEllU5AvVi8tXgD63Cs6Xl9BWr+BOXZV0p7oXw
GI0OOud2X+z/CF2pgvaGQOTutwHHsNMq/6iLR82bFVMQ8tgBf0VcuXk5mhospXb0d9Hq5In1rtQq
Jn4MEroe4NdwO4K58RqH1GrtgYCWI/AT6zhqxCpa50XqSdEOggC/xS0AwirjD9o8bRGr6VXT+Y1e
72+X5YHhVLoFQiTr918XJkP8B32UNAjH57d+Cb1W9Kr/2FkScHoPUKKFS29yQ8f4tLGtk3FvVXsf
aseS+8KkJhl1y58s4qyaZq5jt4R5fnYjvrBIcY2x5PuMdExDnoTfPDku5qAM130aVTXK9SL8ccEq
ed+VrMeiHqod02Trly6871ImKTR6EAHjz4q6i2NwFD1Jg/w+13hhFj3yu3gEalaJMzv9IkF9vwAe
tGReYnggppaZXVfC4meB6XsCA/sKFxobGLF97bXOtH2iM7AIh4vhXaLnnp9lr7IM7rn0WQUDKrWa
F96Njk40joQqpe1OJ65WVk9Z5Zea9oZ+JE9oWs57X2kznlQpoWzqBom4gX3Sd33ZadiljU8zKK6O
uX66hvmSNrVpe9PcXpn0V5umDHFP4F1JOzLRPA4wGDEt5O7RwlyXHMvo5ZHRVIpe8JHaQzrsqtn5
LLdpfTFIduCkOyMrF6FN9e7bvNY9Q0iou/O93ZhjkmLCCtzANJmYqtQ/ld4avH0AdVtoXZjP7MBA
rPFcajrjc2f8rayO8md/Yj/TdW9GCcH4z66eaBLbW7ASfRGXA9TCceHmYa5fBOVfPfZPRzQihQyF
+kZ87rNQcP+fLcQsX1p6b7oMjhNzA/vBmiBzsf7XL+yiFj1N4AiSEHmX9eKGy4JwjFFXfe5tnGNH
S81g+ug=
`protect end_protected
