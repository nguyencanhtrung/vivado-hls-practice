`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
esWyVqSVuMAGJKoS4oHsSvJq+OyHLEFGGtv4yXRTsOiAok/+LCbILT8/Fw845zZPbSV9oZS9rNTJ
87sx2xBiWA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nxZp6klYNJseaWdIuf+u3WBB/P2iClllaDHVcpEV5hWEBWYFK3mizFWvozaTq3htjOidGfYi39h9
W6m956gauWzoGVie9wgmGXQiu0ZRg99OwW4ZQwPyAsggrrp4vVR+HC8zvvAfpcErwOXVHdlN3LxV
1A3I9rBAZp83g8xLQ0Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KwViIstRzVDIH/XdbGFDFjRMSLytbcYHJabneI6aE/rXFAfEcImKeHsT5dblZTJRAivLAxpWCMvn
jifRSJ3vB66VlDr41+4fuKa4YV9NcrYbDH8huiA40/Q8MHxqwZ2iPktqo1YABpKXQDYG2m2CJTgg
/zdPrWvmbYwl0z+64pCD3yft4rJ1C8gDAb07OPX3AsJu7iAukOjyb/PGCQUb3L+JlBFdLo6DipSu
wVx6hdZG5OY6xuwpWNOwKRs4a2jQlo8WO1vcL4Bzt2B618wiuIkdZvOgx2Wmu/3NpVPcYg6tz8Eu
XBCZ6QUDewGuDdPEqIMPIRx3rYpt79anqh3jrQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lavMUGPZQx9gBEQxYgRBD8T5j7X4OgXaLVriZR6N2Gukgtg8oHGBO5uklvW9Hw/LIur1HXjqnFYk
BTg0PmwONMu76YmNPp13XZ7/rE9mf5835uarPH0fQVNHizj+CHqgfj1liTfChGe6XhZDb9N3KzHi
jQ8wPglXIvKscM3DxjY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rwv/DFTe/x4zcKJDtRWJw3MNuYIoulmC5+0DnLoXUAWWwBFIBmUGcdbqr/H+6NzItbguioRHeMDf
wUNfxN0pTtpn9cB7GbbOTtsONf+MWre0KoBIA+E9JPNRn04j0+DtGjZ2g9QOUu20fs2I8WKY6lja
sJAPhA3BzAc/E4S/bMeoPt3+bxwJd3k76jxDVVZUTi34xHF3oaFWMXuC7g+0/cVtWP/X1dd6yzQr
hIDO/yGWaqyxKEzAmm7bWxqv4bbCoffCToOIXQLh/LucfxRiok+ptpZ3WKFJuedd/J+5ZxMRS2V/
yjJac+K2pv98Gv7H4lxqjDVzDTy7Q5Lc9vVaeQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5UIRzMOAfSqdU1i1yCtm69UpbTvNtvk154OFt6NjthsoqdjbRxfws6yaN09Hrk9BmZV2NpmQZMj
zKWCLWdNcbOWZ9kCCsR8EgciGi4y/2yCfkMu09N/dzTT6b+NoFBX16DWyZOvYOi22fbHP0iYiKLB
mc0kPoLciSmAocw13STpVgnCANfB5FRroSDR/tA5rKftYV9Xs2D4bor2wm00N1drceQuQNw5bu3T
OJE0ORhfv9IwRewj+ptYu1sGRGpMaPaCB+50M31OQ8DLdfAQJ/vPLAEILRv6FVEP+Ck+mv0p2unH
FTlbw+c6+JMikg7zF11Ltokmpuv1xRMLux7vQg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7184)
`protect data_block
aqaV19TnAZYd8CSzNFckqCOlODqZEvONkF6K9nGPZsYu/i4EXdvNGE9CqTrslpCiUoE1zzHR494H
b/DYXUoZRAKJd+diVuVJrrHkEIi4HTM5H4s0MOsp2zXuVOn5LZstvr01hD+x1JPounwqHvSzdnsW
t5rwFa682gex9LRmB2+CAR/N4csYd+r/ejYaXEdwpbsBYloKB9HoshheohmWH3tVcXkDJKJCWXi4
XUO0e7G4l1khSgeA/4XnegRBkd9O14vIqJ5aTo1H3nJQ45QbxNJQC8w8ggSy8NuWCmuClHQWCbax
gLRWdJC2ozRExtmjTdF84Usy605/WSzS8eIc+JX8j7PN5w2NDyWwsQHY0YRl8/PIczU1qVeqApnR
+5jF8+UYb3V6IHACsJhIhl/8OFNPJF8aKOczw1qbpEOTFTDfcJ/szpOkH+gsgJVbO0zoWATvMPCN
VzU7WaB45nPuHeh6DowM3KGs9Dog82hK0Vle1HV9ETDyi6oq9wasjju3Qnlk2nuG/iSOzgZZ+SNu
M3ay6kEFHSeX4XH6/4n+d4a3hr3jDd4wsO1cSFrtPdz83XB3XHvwV+LmnI2RIPiZKAHE+k0TSHM0
o5te7Mr/rQklfcCXTfIc39wNCEi0bEuhHbtbKk7r+iTdZpE1O+S14FZk/rKNde24cRyvALEzG3oH
QEOATR5a+GXuWGtLtI5yqfuTsN/iHMbaYfUc6PgEDICFQ2mRxpAMG2qTCAFMjumT/99OvWSjjdZ+
T9wjWOlN189Tt0DuXv1IqpWhRXr87sPCVuQG/rHfo+/XKUespsLLu1jXUmZ08Dcq42TfwqA7DsxH
wwJAvR3ZYFVFxEnXuOhcE5wjIzhfR1wcr2RBoKryaLaEM9/2/vTWSOescA3nd+3lrNowY6lnwWyh
t1GIEF2rmfk4myHk5szsaQ2gr2o/Qzh6QpsbijdmSUxMq3Ah1YtXtNsBm7dsV1ytpv0BK3PeMh6y
oTrT6Qul//L3ICBu/Djd6QVDPaYJAw5mawtez0Y28+lNrg8ch9NFoBO3ss2CtkqGRNyndQUQ/Sv7
bKm7jXCmN0WLSiCg9DEHzHl6/PxCKY9LvBGKHI52vITFEvo0wdoeLoB9WHSMoID/vKgOm4pZOCrb
rpzloxjCp7qreAZPWSpeSIihdLsaMC791EAT5SjJr/m9A1ZbuegsLjU62hxcqt5M62ycSiej2Ufj
o6Yo5LjrdMQIQrai7ciY0yJWg6Ou0jS6u4D2aFk0OfapG1AA5Vlms0thbUbjBg3swxS8CFXAl+BL
usL7vFwA+CI2IQMBfvy+kYHBJcbOn/CZ/dNjCmWdAxs4vgixBI9G5jsq0p+jfLGxIH/UwfDU2xIV
uyBAcAy5/HC18kme7nptHCEaUZ+Tz57n0ldiunXmjUqrBQVfF/80niw1a8ut8LGd/jsmOdkdpCZB
l0mmuOkJ40LNokMXPxR41Pl50Fqc6m6TIeVtrMy+bAOsGg1BG2HHq2uMpq/AOuoLCVhEcVTn9Hxv
N7dRkSapvhPoM8EPQDmnYpgfexcN7U6xZaC3bDOcqHp7zkWDIUhwftmM6Mxekb86048wBJ2PZdH7
jI2tcWwAw6KS2mbDhu1dywv44PtV6iuyIRM2EBCvXWnQLG/ZPXNgLNfSpYLrOIVJXd8dEnAOJRVc
c98Lh4vILIzJaxRdnn93mlczDcUtLPkCpfDZfdWF0TeX0UNVnrMmMON9/yozoimNVM0ggYkoAsHl
DylGWF33S2fsAxjmGIhxxvPnE1DgyXdqEBcTFXFA41nljHr6ODrwd0KMd6RQgHW0fY2VtK5v4j78
xrcqmHZNouC0ravOZjkbWC3qUBIw/+s3aejWe8fCdnLXro6TOShqTkfeyW5Z5dOTAtGg0Q9ZxxBu
AUzdjCWeXdd7SDKREL9pmAZCa7MDWPNNj/7MW8w0c5iz/UHu0Psi/+y86TriTTfoc5qBX9L1YG7O
sKWIO8rSDKZDLtAhUiLYIEt2FOWNUgYAqEFXKEU+dVpXEOmD/VlnyHsLGf4qG50RgU3VyNpF05vl
p7qbM5z+VeV3LOjOn6SjOXhZ99PCuCOoGylwSsHArWHxoP1gZCJx/90lKBWoZBuDg1rzpX/E2ww4
M18ENNjke1D8eMlGNgEHxQEAW0b8HwNxmr1h+uVgyFYS/xldOmQUeMYreThCNjMn/QyHB04dLt5w
q266TVFF260/gTNpa4nKgEBiQZ8IZM2B4DuGPXpkeuM76nd8pRUsqb9EsJ9bd7bpzWWofb7TqHiE
9i6/ZOim8Zk6OEs7qr75uHLod+iz03If/9+dtF7Cv5OH3CBKOniiY334eUr34nKHo5inU+/+12ag
oP3uKYANi3f+8DoubTWb8MpZseCzsGMgTzt1Qr6Linu3PGwWdq+IXUv8vlmGg5eOxr4pwJwuLWnj
hzCrK6SlhRJ5u3gOdGFVKmG+M0a64eFG79uV9qACISQezsPAV6iPwjod/LqBBQFMctkgJysy9J1Q
vpDF/1r7z/8zf9Le4Lrd9m9K8UooVBIq7xofdiGXGTJlsn7K/dV/sUx3s36d4TTcDjF1P4sR6yLS
Uz+w5S5ISmV8szjqB65g5UwN+eeROIrGY8KGC1preEzbqBVQP5V1VQLX2vPK5EmOdwvtW8XZXk7I
jxlhDZiPRVy489hO0HsvrBju95YPRS6cFdTs4IEXqLIt2u6qPocmDQDTmyaHW/okji7DGusM/7ZU
lH0hG7bmbsrqQOYEqKqMgFhoj57n1HNpcdCdG+lrES2rL5HjiHCV4OGqtcqa7rsW8N3uHqQ23Zsg
ZCr6VL2KZYxqQOyfN9xHdbiHI5zYf+ILmP9IZ6MQPl/vOCS4BcJuyEQ1cbXUoEAV/9ErwGFc2Pq7
3q7N0NBZncLTqNzQuJkePLsDkb8+SXIZenM/1k7X0h4WPHstQnBR7wvof7mzz4je5HdVbkIu/J6e
P+OXCXmXhFiJQSF8cL0ge6A1WndB+GzYt7rYmjeWT+D9uc5Be5ct1k6mHWZ2QbbxcAVPd77Qgokv
TCjW1bPwWmwLNauyb+jTq4vBJennNUWRH3Gx68rm+493IDFF+nT5XQMSl2wKzdJZThBTrcyVUMcy
eu5NOJbZSVT1O3pEmw2j/oxib8MX/0WjMwa0mwljbioDDOW6fRUFm+Hj8zs2nPf4TXf+BnRc/1C2
rwpVSsNIc6SwZTdd9zQvDX3MhmDVqzdHgqllSeDe18ggRei2gyBjffSLW/xJmsyOKpkxho1DJ7Lb
2lhEC4nz3ipDMYOHX7UDbhpWnte911Pa7nLebWoQW+JISikSp8x/QJpYOWnOgmLY1Grjj1vKMfX5
XqEuy/3zDtS/UGva9Hy/gdqsyy5JgywPxLhN31mhm2/vOgjKSVmbJYDDGj474edwWY9itmG05qzq
6YEBU+aOfOXPOc4b/bDQi03fjquUl7GhcNH0FiNwecY9CdM2qxvommd4FVRHjUUDp8wkcggH0FOU
3LxmCxOmeny74GhXkI9EyGYZO93QI+loBY4G//3p1LuSuiHLUKH7baO+fjc6ir7gpnzGEuXSYIa2
Q7ffwIY0O6SIzDS3yQl2kcEQBCk6UwkzI1HZRiQtZ0jkjFNJ/ojQqAr+ai5Wg1/PCzbqMTo1OpCD
yA492Vh+iQ8eKlqCCtrWkQl7nz+nG5ixZCzp4J1WilV/jN2R5s95OKmMOpc3BlcdNHaWIiXRViKH
du++FhCkQnduV+9V1RT37FbX7y7YTjo9MFvFeLmYkiAqzlaxRi+7WJTpa1IFxFxZ0MljjqlmMmi3
zY4r2hPXm7HoLF0vEsvrK2y+BdpB02YpjcGIWUq29yDI4EN/87riNXr8beThqNq+n+FXWSY2gCsz
xot4zUUzi8XhQtJ9Xppv56mVyqOLU5epSl3XGlFQIgURsA+TPesxskry/oR+8alDD4IjBPf3vBb4
hi+tHaxHjoQXotu/L5fiJs7GUwD31Xe8zmQDkSqVVMQPc2+K9yF0jc/oWm1VN2n6ccI71IcMAZYB
8fQnevJ/v7JLLMEePr4poj2421w1XkhkhS7cUOdrRfk5SjyjKYa3uyEJiraOO766fApdvHJO+LsK
N1c9/STHrCxElB+IQrqNFIEKUO2cad41qvmv+aUQq98wZkceDIcAW55+5PCLBZXrCon6KK0lwl9Y
uarTlWYdlGsdYC0GGQoFwB8ua8Pvz0tH05wK7nQsb9E9P4y2/dGHywQZoOGQr9kahLeV0f7mE2iG
nVKNlYlhFhV+TFpd5s9G24i1asKqgzb/hQLdyysJ9ReF5FVCIv5SXN00G1LWcFaVM912YgM7C7ju
jJPWjxjw0ZFoI5w+24oQtvfDH1PCqNyL2QVujQ6FZLucbau+dgo5XNY6Oy6cydAZFXHKuw479VP8
99vfItiv0aG2J+RxyJrLQAPb4o2oA2qm9Hlu/O/Uj+Z1B2XprvBdINKBssOlHGl7a8VfHsLym8HF
oVVM36pB3HToEfizdXJgMRQAnWxAibHeDPbPEC/9CFdD5hCKIvaajzpf+x/1X7u9r+YrMLnhEloj
g2lSoc7TXSnNecEdtOfGhMJQWqroN52GUkB+PO7kN9rPFoJL1/60toiF68IMQbcP81XKQUBx3+iu
RDK8+v6TsQryPOQsaujrYLDuWAhoq7H3K73B041J32sgHIvzZVBM8npw7dwAwt9Wae3BoN2Z93Ra
W8TdgX5nRjZM89Mpws+EdxX0fAPAEvJCFg1E+Yd7Ck9EF9A6rmwx8gqTMG+VTu9KhmWDgIVpHsdL
Fthkd7dKgVu1StB33XcPhzJYnloO/h9x9UyxSeYyxD+h5kRDEWDmT6c067LljHJ/Dx/VdoaDvhFe
rc1vnX7GodPLgBUngk3LF39VqYlAcGAPNayVMt6z8iAxXf+AgcCMYcGk1A3n/J37/xXGj3RHu+03
mSEZZfArOYhDh00NXLfOkeGCp0TzRwhPyUQAt8/NXqbXNYXZzSwyMsDoojPc6re7nVQ/11EuUwsI
KNd3FXo0Rc7FqDqnggLUrw6i+uEyLu0L9vI1DcKkEKf86mkUo4VXmktGadqhu28z1VFSv4y6kUEi
WbO9Ti2xZQyAJodqG7VV/61LRzBF9Bt5/9tfas7LgENxjhfgkQ4C0qxWqfuFNc654tTvoUyaCMY8
4NQ4p5dRvqQn9gAlsg/uyuxAa2b4x+3FaCVTlDfqKIq8aS+Me20/krK6LobPwm47q39+lTesq4uO
hhz4yr9BtJDkzQ48lnuR0oT8sxLWnS++TxosZi0cHOR8MGpGcprnSbjHdYTaX0fsLAXJ1Yy1Ba2D
fyNVxxVhm/C4JSqJC+VlSI35xKxx2PIx5zO1XkuTZUjJP5YSr6fszN9tDDY3VoQN5YxWG430li+K
1GFo8wGqy/EkZXhWZ/ftPHYi11pORte6nVitLtZ0udLXg4YN/lLPaPletw2ps/cyPD1INrA7iQla
cgHlI/NgTLrJn7/PyxtO3yOzl0km5tvKJKdKw3welodFxrxH7s+LGSo5AoLwXV7Pm+g5jltNv3CX
QrX8YmFEtHmhOXSk/X+th8HJsYnO8m6m6e7QeVrQOA5n5ZfNdGCDetQ/R5nrVBUoXFVe18urF3jX
tmFu2KjmoP8j5dO9Hmm9JAFmSFuUBqLvO5bTpkkxV+5tOZmC8fPIjz8yPvJZ9w1fjApV2wYjCFYz
PtTYy4piSEMG+mppy4enQjFWaC7FTv0dz79VvcNZLZlpOGFO5XsFZ4G4o1o/BnGc1JD6qfvaaRED
vKlEjKhXmXQcokFsZzy+O0n9lMMCs5b9CZ266g+Y+Jg5iHqEgewi8XjQOPLsUqltaWBEloYeT6dD
08ZVvZRBw68el5Ll2SI0YAz16ao5dfAa3WRxybZCxsOZdvQTTeKor0whsvVl6MgTcgSHlRLQPST4
SCeOTb2723mmbkGKAsHV0G/9KIRG/lCENAicWVAio+9n8WEI5lzoDoOJGVOGaAQv5jbEQY+b8wQf
YA0U8qwiT/KJZctxOEunyTQmcnI5efOqYy5GqVUTuOn8G8Jtbpd9uucBJx81Rym6EIJxuYVETF42
jigjL8GNiRBVVicbGTAgmlDkmHSljWOTjqOVFKGOQ02i8Jw6n+LEQrMQ38puLLwaMn5hlz4x0uWk
ohCiSnrBdZrLRBsWxOh7q69MSBu3hHAUGhz/2tUC5mBeC3sq0y5HnlTqzDxR5PGkfYSfcaym9zFt
ak6NDBO06fV0FHC0AgTJ+1n9Dz7eOfwq/Oi5+LpGuEP8EjkyCdtL0+St9SJ3Gu6ZbILKfdX4ILWM
PFDzKuiKDuGbj+nbO20sby/1zGS/+Ln3XDW73EEnPrHStQ8wNTDQLMzyZwHqpvfErfrOUprvazUK
gyN6N0wUE2NC4kVhFFI+K8qSn9optnBajY7H5rmC/gxJZIKUtFvELaSi/hiZZc4P3CNiRCNfgBcg
gQ3fk7I/IAdQHz9SsBVUUAsFJDaqKipfbeDTSlnWGifc67LfyOM9KFl8x1Gw5mC1VZY+vSU+bnBc
IzcrXEdz34fxQvOOlkBMr3NQaufB4/vJx1M5LS1H2tS/MvKjrQMpFGD4dqPQ6Pgv3rIQsdYXSxF3
j4jX6RdcbNFsPrEMWlcNdMMNBAsa5lG8ebpoM74Lf+IpjhvI6tUG0f34ssKvV4CoQpB6RsoVv5J8
13b5B4N0GN6oUAyeQsZJJvpCmbDxmieu/uKAbzymUQgUJfSuaetDeg6snASZEVae4zanVXG9exu9
hcLQks7+NbujfCVeRrnc6i8oJgiI8SujSHa7gBjNsCr8biyftp31V876pb4VFJNK/Y7WT82hu6Rx
BortBqwiBi0wQnfilrzNUOUjz+E/qFeYH86hHaOwdN8H+OrcLai6Jz6lKJKJeKdWlulvPypyMIT2
dncN+aEPuqGJFPIoXAumxHiY4FizFAOTnukxiDoekQmOseMbrBQ4aRod0jl+BcaFSiSl+X0/jCk4
QR+2TRDsYzfy4e8C4bas1dOKLBvH1tPZhKxhRlPpKkOGLe4sSRYoE/rGnccmG0t7UaxTr8o5OPfZ
8jNtpLp5oueQHfbAEZZOUAuqYRpWDLw3vK85Tr0jI0BOxOxe3yqyGZ5kf23LGS3F1+cyQr/0vPNi
htFuyu/zb5vwpO4bGgFs3ViutK7pqeCa6JN2OUGYcxNPS5zYYEJFMDzlPw22DwJGjsRx6keG9Kmu
KBfLPOGraavH1vwFqiBfOoHisk9DDFdzZ568CYTrk1zZRr8U+WdWR2k7UGrZJ/HbGHL3WJqpMwc4
xlUxr7114k4fW/1sQC8ZVl45vxNrH7ai0MTYe8sNQf0GUW3gprns9Cu5Y9qFykbe0BJE5zmFTjMN
hZwX1ILA27QOUYocyqNqe1h3eBMxWs967Wy0UmHojv6qJMwVfuY/hrR+PyPeGRLpiUXlu+YmzHTe
2P4MYcQ4WsZx+BN8/p4REvaCQ2yLfNxL73a2q0UljpyjGlLoXrKr6vMdzSBEKFMegQCAOl4ekA4k
tgsVUswPfKQB6z2y3il1+At98wHP96XxKc2hhtWDSpUdH6S/7xyHVNfj+wikmjf+P07rniKhLJb2
4R3VjSuMhT9yKxKEneVylNmju7OmQAoalhixdL77S2inKHqEhnJf4exT8KcrYc3LtbeFoZqv8d6B
+PO7R+OpMzcLmH6dIkxMQtOhgLE7nzSskNzr1p0uY0U9m9VfWur899xuCpW0wCF/d/ky8MiQ8Yk5
SiWqfza8vjx0CUvEF53+57XOX2ofPVHVOLSvz/5kZ7Ya/bbmD1y77yO3dTXCzrpfPIAtNX6kfmCz
xxcVf3Qt8kQf01lRMCza6Kethid9C1kjlTAJwch5D3FqsBMZ9XpMLREKlMbFksMKUIFOoL/vdgtN
CHGMlvUXMcrnY+tNVdoW0X4TRI8MwQDE9S2J6A5OhwXyWZxVQUg5S2ypQ8D2RBufkDTBEBT/xtbH
lbqdZ/fvV6dsKKxyefWTMqItEgjtoZ0i1ONq059QHgmD7X6RbMkgGtf0L0tu9aAsuP42heWj/nQc
KjX8GQhufiQK+p1PYEBS5HeTZlTrZItUr4dLVIIIvaZk3VZQjs4bY4NuKVEUGm86aYH9SK0vMHq0
065KR4mPP797T/j/q5StxFyKnWkiM0ml2H3fvoh0N4FaW3gmqFjubQhg67nnCD5TGtTxjiyCoyrs
4s5BG2+Q5HF9qr3Qk3d63fo9efGyVGOL+ixB3hQey/v8ifP6xpX9TZ+AtoU9JD+SypB0EiTzWnA7
vDRTELV5ypZFmqxfx6oCXDs1y5nxvFkwgiSKcKjGdVhfQo73pn1fYWkvixwoGKqjw1b1WGaeSReR
26VLJfXRQ2v5KY4o5Ho6KmOgO3GLeK9/ghHTC/pLaPqb/D9tW3qtT2XWowRW8bLMqg0I4DUieiVW
WIEK9wZdsbVjWjOtIpMc6mimIdxHtvidzB1rAcLm3jPjpwddZJQmE0wnHLcwspLrZYjQ/uauruv9
a/+WZuGrBIhafZTST7usjaS1Y4zxqbPvEjvMW6IArrJVwdDf0Y0i1Mz46Lv1TiMIpAGjgp5f76Yu
zmjmMaJxtcqQ2eSpJnHcqnZ/GYpY9CBfNiUR4PE+3OrIvJc6R0+cBGBQ5MFguUzVSbq6ymDFdozr
ukTLcSONt7TibxD39dI+peMGJr8cd77whEiTOjzMPXbUS0LK6ygBY2JrPWf0NJn0bY98Ms6GAS7d
XM6Dn+IVDfIf7X+NFbpD926s1EcVnmV11rHlCmDaQZb6T4GDS+Lmnkm34sqH1J/zQ0kXgOYzSd+L
6Pnuq8tb0azS6mwAxKokjejnVEbaHb+8k8Uae9n9TJakcWvT48PdypfDdyteR9D3cIjFnL+bLBFB
mPqZ9wTP2yaP5CmWchuHoEYhczVAYwWItoA7pj4Pa2yfBlDZGa6ekDes+jO83e+xL4jnvvDLdw8m
Y7QROYl6cyX8jM570zJk4g0ZzTC66NhHBEZCPNoUCOkGEizR1M9q5xj+G/dX/bhJ+ke/ozND6P9D
oYfw169WLNZrkdrGsB+esY31h+ZcCxIUM8MKEGxHuTWlc+izWSPuuXSBjIxGrORI6+/voekMrtg8
7iZXjfzKJ7vC9jyrLgVq2/Vx+FpHoZU4NJY1bK5sj1mGMw4zHx+ntii3iNeFA90ykBUOcM9jcSK/
bclpIGgqyDsT1KDQ1egQzljrCs37j2quevYK57zqkoV6zdQPBJ7qeYyMJY8TjO/syKmoln0UUgz+
SPBx8Kdd8NTjHvKv9cBKITTGpmlwv1J5tlMtEwYX+wx4p3Cb/tV7sDwFkI13Y4FjekhkKV5wklzO
jSDopaERs7II/Z3gm6b8Dqs/y45yn38W7jEqSy6ZZ/yg7zlvAFuZdc7opqAnPJp+6NglynSX+3CE
dJcRDxLhhumnbwtUM7N06BNt73jFZGP9rZWJwqSVpXUBge9rowgCtPLTDX+9dTQmqd5hwfFuuQd3
Hrnptx04+IW5Aypa/6qNFy46EFy11k+cyNyQeIRgMiAtEeGc/aNM9h/rI8XDebmoHsY18ff+R5DN
u04=
`protect end_protected
