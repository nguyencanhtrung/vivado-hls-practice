`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Mg6xSA+dlOFbHxne1ZshpwlqADvRNdfnP0QyUcfq1GAwHMclqGC4mrKdlawRjzK41rYv6AHRAnIU
RBONU8e9CQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hXBv8p3a+t8pC16ezuhif/vvO/j8JjwzgA42J5TlEKNuxyQxrbHed4Y2tB3VbGrLUDoc8rx/jCwy
9QHvZYNqUqcE/8XgRjJEr9/cX7Cxxy/k5bjtcn0hfY9padivE77AA7kY8DithSOsBPi+MiDJBTFG
L18D7zdHFg/OKDyJeKc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JV+KlCuuxwz+SydG4Z+SsYW8IXTEkav0v/Mbx9Y5r9wd6uaIslo1zb+zIB+eDuk72bKaWiunkGWa
CSfr12yPAoIuA0wfr1FqC9+Hq/un8BDaNmKh9HK/5hkWZ5pyo+40PsGMYc3qhU0vCMTTd5qeNToI
7ScZ47s8K3i+79yHxpWTZo5bOuRKfznI7bE8r3k5i8+g496Ess14vw73tvE1+znT+5CUR4OfMLnY
PX5TBaZUhn8h3P1Yf0N4iJziAMjARzFz2lwyBLq8CEcAGtFmMxDNowdKibAOOppBBM7m8Hk1i6W5
loxekm6yma/e/UeZImZ63RRh4vSdWOFYGiHOnA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vyU3gdWtAFyC0iWQwvtfCNcUkiMgPg2yyAMqAX+j7TYeIWrvqta370KSeEsX81T2j4mByKB+u9gy
Gpo/iUJx8gJ4RguADq7tTyEQAln8RM28GrOn7DZRqxavojrF/RE6AAwdKHtm/7arWXdK9ApL7Rml
tvDe2zhXmhf8ec0supE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dSyiGob3Yzx6m4tkM7k64lW8GyGniR9t/fVEti1tn/EUimSnpNi5EexU6HM63h18TSTH++cZnKG3
gw+11tUpOWofWz0TpVFc6hUKU3lFF8N8f/yjE7FFXa2Bly0CPC3EbVNMOI325XonAX5tYgS2WshB
To44gtnN2afSvV2o2Yv7IEvkrOWZ4kTQ0IxePMCrTOLIQ1LGySyLye5oIUM6Yzek25VupM5LsWbm
4WIEB3K1O9tRKZSi6iBWtsz4mBFn19nbwSGC9CiqqyHtgmbqx/1/+mbKSJpoz2j9x8/n1aWhySWs
02yCkkrp2XRVjidKvujtxa9MNTc0lTJ8OYd/4A==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kbx7ytl+MrBv/yhvTT5cEeggzTJXOaPbZKR3DXk43NYTg8WTbsm2b5K1oGPeR+/iYcL8N6INW4ur
aQI38gLK8qwxFUxbGCzp4l/KtFy+JthH0b6MvtpdcxSZHSdb1oBh//KGCA7geBzjp+MQ7OWK7hLx
Y79R3SIJihykpEZiQU063pxcQWMF3xN+g1iBKnEBp4ykhDOE71DTAt2L6A2ZD05635hnPNoEXtdz
wl/iE6tWA0FSixoCCih3hKcopq2Nxt+7F+71iHZT6J5Kvpz2pfluv5qZM9JEeWqp1PyuaznSlBVt
35nGa2cR7alvaHSFX2cNXMJCyZ51SJhjuk7POA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 168544)
`protect data_block
J2BX/9ZMF155YVaz1MV/oRdd1+x7t1OL05wHtka0dHURmW/W2Rx5PFVpAktYd6ORY1VFkZ7KGPL4
BYs79K8SstQfLTkhrLS1fVixAuKznAJswtOUmYXjtlGEsB1P2Mb1+84b/Z99+979yHolmhByVZh/
4CjHogkSqVOYHb+a1xJ+2DE21u+eKiGoHtUXpqVgTWvspWTRLM71X7EijSx2cC7Plj6vO+f9ziJy
fVZ2h6mkR1n0o0yAXVi5HnpNmUpwmdR2QU9zJ7UX3+1trIR4/tyBMIody5SvkAwNymmWVVvohuKW
EiS+8Z2v/tHMS3gjl+rXZqeOvDgnOJmPFJy1yDpqvQW/hwFSrmsxF0qIRRowSzXnC5AUw8iPvrse
GkNTzK1CGhciBETX4QcqBKZSopCqDrfxqcM3vAOpkClxgZBB+g+I8YCH86fzidnwP2amZeDt1QE2
IrNv05oH3yUa4FY2gk9Jk+rP7uQ/pAv7Oaq0BtOFDTGLciGn1Dn3iJEa6qBh0jcpcIYWh2AeHPUM
Q3j8Cgz3izve+CIEryMoEMJsChrZOYhXxvqdOrCkpt6yE/U0ed5msXRiDzwP9+YXU/C+Qjue6M1M
V1LwBr6lNhxhkNDk830jaXSGRzueQ1IWzQX6+2V98joxNpdMC9kjkaEsr2fG7PgeicJyCUlYTg5U
x8Peuv6s1cotmTypxWHlW69V3y3iQVyrNe8jrnJCUdgzwQoDmwyJ/AoQoajPyvfDZW5EAkh2ZgL5
0GAjnI1860MMyT86/6Tr9DGieyPjeCsK6aKMYgSYvWVzcVGnYedbEAuPkvaNKq6tiSehxiv9xaNa
eY5XqhEidhb/5tmFoN1uV5zAk/k7wApXXcW50ykj8Sggz6Mim6+IgUrOyuoaD1JWh4y4qstlHQgW
YKDbzJWbiEctiXzSsrHtpa57pUK2WTOSQfS/cT6/URTLCdUz41FQTvtzbC2RIoWJLwJWK2mnDlui
f+6Frt8MogOhgjUXQBnV28JllPclkS1cPTXVql312CgKptvmy+QSwjbXlVOvBwR+ljNwz0R6gfD+
0n+VwgUG3UGD/D7f2IvO+ViZ+egXPmxYEyC06Z0sRuG38ub6za7Fcwrgusg4jaglx4+k8Ngdqzmk
L+BtekWIYVD0uPewqODD2i11xAtMSvCS52SQiLbqbe+vVdd5Ukuv9bqjAsiaeX1h+4CzR7kkqbR0
aU8DZN3bzUCweo9qfCkXbkCweSD/9UvyBrlhNDuCJ7TOU6e6r78zvzBtEHgmhYYr8gapCvVyGplS
xAgMN12kVu/NmTrCfJ+ClNuvBACRKRXpSM5cHnPHHldolXZXmxEQQrGpKPwe21OPiDvJfybPy57J
sxRw0jZPekK4+dd+x3nl5CIw0TYsC1b2MG3t8/FHyAxJZjD03fPUNh7y6LyuzslWhQA89LguSm3z
Pougujv5Gw9phMYqkEQa6JygivWdr+qs4FPk7C/TAf1ztGqBjzQXKTw6Bs4cVuTzCME87hHEbFS6
J/DG7csT6o6sxl5g1kQ2q3rREvjyrRuFAgfl0YJBRyw+MnjzT7fqCph1C4VywFJH1HJNVzmdgSpw
LSMjie6z9b/LyEiYRyr8GBE6nvuQNazZvOSalgyzQDMCi+kN1cS40K/hA1QDj/IgHglGbz6LwvjP
iJ/7/z8wa75vcPLKXNYj7hDHxVRUWMasT4txuhTScMzumFm3tXg1Ck9gu6I6J6HJzKRDpAGDqduB
R6DgdQkdkOtGOxmSmLsPNApfL3NQpcf61eQYt32g2tWpeR4Krhl10gdBybzPcHENDsY+EjlADDf7
Dt71/57xDuUwuHRbk5Kci4G2rPxdfFm0koRPD3b8rTHivBpE5UPrkEj1vOvF/ciTTdYjJbx6nUBI
h85Xtu/68C+Naq8g1AINgDRd8+ik6PJ3c+I/VF2r8nxuBKZTqacAQs54hxeQqvzkmT2p2qI27AOf
tOdxniETicY3K7LRcFq80YQKyY7k93VVjkB0qHWpwqQCxLFMR+QZdfTxq5QRaf6IRCyZso8WNfLV
6KQmyPiedvPDUG4EwGEwvWZiFSwMNbZvHaWt+j2HwOI1ca2peMVzlTTSdaDLKdcHxioXPZlscoAL
F/uCwp2kYXfIL/vFlxwl58PvIs85NUyRi+96WDP21Vn3zlYLDwO46D7FUEyn7K+yGMIHoNYWc7q4
MoS3i001QOwcDWYUODXl7GZhnbW7+tqdzolnk7ebNLACZJK3ztnrcbcfeLwpvEmWUH+tAAqby86J
DCp0Sp9nxTVeCtytOQSIHzsxWv0TDySHcp0L55u3i0tnrDtc78Pb/VFUkdBAB+sbQzGgRwG5qEeN
pLlpo8XGx4PtflqRk0zuzpM3Q8tgOoO7Vi+ohlCI+N9u1HRsEIGmBKjp8q5l5yjsa+3Q0YQa9mJt
cdmjbUVol8zjj2Bo6HmyYREBsnX7Hue5ExZS0AO1ccPKzgjEzWPrxGTPZ1lbdmO7pu9GXWMe6VVP
Re6VfcM/uvoA37UK6jGgk9686Kxt1yBt39o+76Gtie/EXA+I1YlUnvcUyN0JgzAnM5/i/2IIgWuy
oLIu4S2Ou8x5GgOD/OBiSYWkc/80VVsPDqhfSd1kuLCyPrNYp5Klkuv7JjQ2Nj9/KBju2hdQ16Pm
Qdi3A/kjsVrexHZiUDhiFJVng/VljMCIR7N5zYn60+nKda1JI+aYxXHx692Zp3eFd6zBkGOcF6HR
cuZstsnvhpBx7D8YPpaH+BdNERibduiBJpdlLuotAKAl+vVV4TmE9HHywotLeKYwOdwWxPr6Rbfb
XlPmv/mtp5cvNLAz7I9FQaV8Jxl85cJmvORSx0f8LQUySbh94CoWDXLU3slVXTZdlAmU6NEALqhn
UuobK16W0fogWlY/KyQEvRAUXdEnJQiH7D1lD/cp3fEf8YI1cu42pys22w/bPr9YAcgmuKnjfgqk
JNJg1rsnN4np4rV+zX1mKACRaPV5rBEU2E+rXM7GoOtBD9dT1MEgb9Vr2nREOGQYyjPd01vfYID4
FbF8WkbYbJ7BKNwqYKOHrDy2yk0fskaRi0wuXlSaCpGXiVNOP9IefqOVAVu66ZcBvl5CXFyrJ+el
J7w1uG5vvHrVKXGdKMZKXT+l5S7u6c5pDz871FnEERnzNFjWUFFwdwxq039AjXkE3h+O0T8hv8c0
qF4QxS40QKATiSRRKDXWcZHGIbbkk5lEPhQauJQjMPhFmE/PzSanuJSKzRFLa56BIeX+RVR1VnOG
p6IeDCzZ+JIpW8nDKrONG4H14WxeqmyVapbyZFUiofhn9Jujli6Gx3kqrHu9YmZVpeEMoH5rZGzR
yeo2vUIXq944vOAxZ5f4Aj4i9DJfeBcFVL4ozsqNW1iz1cJk85C+yzplqWf7hWUZFHTUwUwh4BvR
TV3WuatXqn8YBl498QBQjAKE2btbBPIK9WUkD5jiEjkeVqx3rp4+dAMESr0dM1vy/O2oXgB1+q39
fctrPG1YqIPzYz83VlJcIjVSrw2Ne/PAHbMMZAIM7BRfysjIzJM+8B8mjR77p3YSrbt0SUQWIV7Q
e9o2xOHvIyBQK0hyNr9pvWW+fX28HC2Z73EKT+QVugD3sISVcSutUojSr83qRYuykXRL56OaFh6m
TXQ4IjhvH1gKm0R6YVLkXMNE1iN0Y1oTUHu9x/lais1lJy/hrOAGDs9rpUKajJG7a8KN7AoCKWG+
UHkK7qKmjEsQBSD2oOOhy/ijM1vSzbYp5xH2h+OXQN2WaNQuonAsOSv/gjJ0+bGHUhoVRsgI8MO+
eGyqqVF+/rBk8f8KZKExpgmzFufnBLIsjl+vtgMD2gB16q7iJeW3wb+x1ZIEAzJqE+6pK7yH4kbp
OI7SXNFgRZUI7NPe/Ny38slr30l2pp3uf9a8D2+uiLFy+dSxeiTw5HMKRuIHq0Ve92uO7QD1ldPV
MoYB0cZGseD41hhcTh9ng9AY/p9yIW427y10NyaZAtOU1+ks5D/AIZj18Kerj5PzNnWNsigWntSu
fET0Hj6+0yUGV4GBqE7iXReVDcyWkCeuIdiB6f/dvNbCjlEl9J4dNuk67Zb6VjMdxq1SkPAtqZFP
5MxTLNMmhKqCXqM7x12DoT0dkb3wPnaOwjQas8s7pYdtjQX3kBCubCiDlRxov22svbFq9oPNBDNE
90woeSJphBqOnRYaVrD+3OQTymaFlx1igs/F23DhEosdqjB+Cm89GAQKES4moMidx16mGW0p9k6d
X0thmokDpki/SnXAn5UZI0hjOInqA32IH/hyvZGPwuaoUqjnIIFb9MIY3CvWqzVfwW9o8KtvpF4T
yvm9eVLDSGJ5JsqK2J7CKgCN5J74CuivtuTGVM8ouSAyOw5w6ev0r/nPQ/nkL8+9UsCNfpp7Re7a
x3lhnlliW0GIR7Xnis1qR7tVPXYQVveCQfgaQe9WA75aBbngwqyR3Iu1gtZU/VL6xRmDYwgbmHhf
ngNzmiquqAoAixOV+gibU0ZC6vBLs4qY6cMUGbryQX3dhrksL2tql65w5tKhVG6bGkcQsXftFcOi
j0GIVQNi+z7hbU9WWp1fktnn1qI2kbrte6kH4CW+GzH3f7s4WfJPqjz9tqeuJG9xrLYuiJnF1Bz7
E4SCryy2dBPKgxgeVvRoUnfQdS2hF114jEtakMTMTD2huwebA1TX3WlTBeYkxvIUfC8AwNmotGY6
9Vx5fa7lYMmewiFy6UQJwBMF3ju4/WpG8+PGQ6j8XpGAuyKDcI6b1QA6zeRm8KiuEIL1S213oPBu
4oOtvDYrd7zPeQxH0uwNLblJYTR0K8K0A8QJxtQPlEKolSVMwIbwd5W8um9avQHDw4+MOZKhDcg5
SiTrZ0rd7Hnvb9x7ZdKmcdgvieLWHFFs3U0FrWrYhQkISqywaSRBQmYvQs5fdlLSQ4o8ITHfoHbp
Idal3RL5vMEEDvpiqpGiNouLjYLWCyT5z6/LwhHBo9PzP4uQ2XiaW+UE6Aqarspw8mB7KjmuSAjN
D/v0MtZk/lMSAXG+NrSvoTqIVtmuqGoBNhp9BhZpjnu5zNwF8L/ieocjnbd4CMYS9s/HpanhmnYU
VZYUIkxed26t5Rgv1rSfgAIJ14wQJbI78rFFGz0Lk0ARzrJ+AARTUVEgk2TQyBKyisoEGKU53QOb
bsUQxr2LgiZIxfs14OgZy8RKh9LjLBNdMGG5j2l8sxGNNMZX1rdkdIR1e8oGglbeTsN2eMk9GYak
r2na+T8IiEG2t9a2BjFZRUT67Gyou8uyxhYaq86nfgLYfnUKi0M2x0WxgSjs2AnjmShRAWzVJZjS
zPv8IePCC4Wjca5OVPVQcPt9ALhz51MepOEC74x8CnoM7UIi1zBZRWG1Fdrb5nqFPRmqIwQNkVxx
FZ/tDT/WLhCnROQC7NRzQeRFxlRib/OENg4OxlQCa9aB+3uVquf6XifuCBVqGmRYrXB8I8ztSYNt
qbyMTsPMPq1WpAROS862Pruk6UuBrKJavLM3QdjsjZcbD4RC+N6C/+F7WGEgHzWWFqd7HxexyKIO
nuMDEMGuxYRrkcOuQXFQGOrv10d7l0dTQ9bzmb9aoZG7J66STgvyNc9EpoMbZMMOvqTWHVw/SQ/p
eRrsW29FmxTSpvnao/2kX/WP32B6Pke0iCq+LnhEEexBk2SiJWt1aaUF+dFCCrzrkyOlQL/0yc57
mNk5To6nt7SkncyC63K2nMlF4VOwoFkg3TB1OCnaKgeqYDz+ZXcyTklFBBHqQ7wX7gq92muVOW2k
PVihTHJoMKyDMCboqAM/uD7/xbk2avBgFJT0lv4US1RTqFKrBPSgfyGcDGgxBmzW/SGAYyK+iTMq
1pCNiEwlCWQOJMIkqTD0Xfix0nAxJToMu/9YolG6VyWEe5PD46Qy52WBMVmm0egpVTagYXo63w4X
z6MfEeu7nV26dxvtYfz+QciIOOROqAYyj4hO2iPYh2R1+ZPRufF72/A4ej5wxvgzV1wqh3kyH+f6
VWQKcM2T1LTZOY16aksJT9npWd5zu0aF12WsOj/0WgLlQM0l/A744Ekfue4+r6lKE7NfSqRTlwU1
meWMZVYGTjElYfsUIzEcVdD3AV2O2KkeSoM6vtJMEWwnCu6gETeeuotMOyo+X55W5GTo1xzbQesL
a4pSYA5m/b5mvumko3PLZecBBIkK6GbBWlne//eH/+8eKAhxGg+AyC+a0NrmID3VxDzdyIq9JUM/
veSfwbqb5762VKV1724BCNfaD4dQen5FvE/ihZlXPdYn4toRECbiVn1UT5E91hIazcgsc2jvHy1Z
TzgmxRx1J8P6A6m7U7mTsZZRv08FJDLyJIcm4Ayywmbi75h+8qMobeIqYQPvrGlyDvlqIb5GwUmM
NZY6XLkkv4UpsN2/PzmB2/RhEGKgLeAlGjRdwGENtpDfpDgYCMrXtY2hIhVMTouPq29fwDDlr9P9
/UxD6ZuiAKBJrf1wHrOiel/pWzheOj5Q7WgvhCubOK7fnO81WiFzN0Gdt15OlvHTOZsDMuqRx3bZ
/8FxGrp/VrFJJlxynezwlD2zhD2QLRrk+vqPrWVnlvYeI7bSS6qBywr+sfmGtZN4YElX23TyPv8h
k4fQ6UMqugmKzBXRuLo6FsqDeLn0on02h/1F3AHXVEXc8E7czHlkvDSgUUEgz2E9qA4qqkVdrFw+
bjZ0iSPMOTHAXB2Qyfg3nrwhWBSWJaIGaCFwJT0MhSzG/etD6AX10pXONzjgbm4kuN/pfob81z/W
XuxRHmxCOULMb4U5lzdNtOPttXVjVMQAkhscXAZnj+hBr+bkdMR5QxI0ps0Iya7/tKMHO1cRtwYQ
iUqEBp5EbVI9TWbzkjuOK/I6RP754LeDnTzQmAkuaFtlYSiogakYtfhnJlPUcWh6RIHjYj2EXub3
pZJ/Q5Ywgcs0PHf+glkRI0fRh4rjhh5aRZHEaDaLRY/CgLNJA38URkWYrj7kijA7otFzaoWyH18+
M6THmhy1VEOxnFkWXGrZNzMLLb3M8w9dal4MPGlAOHd/3vrapjVTyOnOSB1fabTGFSmlMZi9hDJP
O5+NaKgAuZhXC1TYT/CrsKY06cdiqLIFcOc/3yTfp6eWt2CfrlWV/IjxJwADL4TsMis/L5/+mDh2
+WDtHUpXrvI/PvDKfT93xEeUEAXe78gV65GLUexb4/fvUFKEIDd7CdT1d0z8LryTQ+o/B+K/amGC
kWyiNndXsO89AsrNFBr6bgATH0rckQ5w0HHWn1u9JfiWwHb83tJmnjdyrSbr3m5Y+ngjyh3wqa0o
zcDfq2fIeUw3ImYU0EJjZPBHAg5WUB3WyzwrfO1nWNwrfmxJWEmzQ/yQEhsvZGkG+Lhn1EXn/jRr
jUJOG5dUoqHQmmVTCIDANHzy7FZ0/Cc71gkWVdurEDb3yYNpIMzGmG+rbrSId/Cw1wJ+R8railqA
3O6ITwTpXNuekEmTxQyXFt8eOa3B83YGFZCD+RQKWih2cY8Bkng0Kh5jR1bMvm9+T5yi3GC/HyWN
79YRl7n6qvzv8FndupXQytd5jtLkGEDNYj48ns9lQtnaUl09MvpWn3wiSLUasLWvLlqaJGLhX+ur
MyctNYEZ3WIqv5Ewvnu6ArO+7scOVVIzq0OYyzdonhQSxNC25TkT86w9ha1nn/VEs21Cj1cURM+F
KsQ3SyhfyA2nOiN/mpPkI5NLaTmf/EKt7bdjNw2xLY/wRNDGz3syJJJ3l22jbOLXmDZtDsjkECS2
FBOwrJNrI6z+yAWdCTkV6utlBp2keIso6Jvnv5oHR64Sjd6z9nieLdHh34DZYG4C2HZfUQkFsrNb
zwd5gvE0M2sBwRYuoluT8pQoIfBgc+EyQSRFV7UEDYeAXzjRJTg7ji7QOtxYqUM7DhSt6KsyyOiW
pRHljDo8CA04KvJq32tDAsY8B+wzsMcbzPE2X4VIZ4Zz6FnrGFfvYZoBaoc4XP2lZCoGLSgsWrwe
zq2tkUeisq3BTA2rvBxjA5wvpMaGZR5Ik89VfnEtpvNyLHqKPwOwuecN00YzcKe3aROmQ2LGhH3S
0YpHDM53J9dekg8SYcEYENM67kgrZbsdlA/sLDMrNny100oxmc9UqnAi5+KnlsWDI/x3oyrLSoiD
Ra0QrYsIdyavYzEcSC3gLiRpUJrN2tl9oQHYo9w5xl3NMlgqIJC+E5Lu7qzic8VV1Q8HI4QZrjzI
a8lXMe/s3e6xq7VW56ZnttdCXhMKUqVYsp+OWNHWM9LvdVcMuvvUa7J9alsYUR3TWaOC8IDHaWzq
zAoGjdjbdNBxNK40kOiP0ktMPT+T98QewVlDngvdCnm1++mx2Ua1KBhrM7C4z5IIOfMIpdLE9S0F
FM2vK87IVsXr8KM3IfUUF8+57greWCiJJecODbnTEPDTU1mngi5Ramudou22WLmrWY3Vd6VAYdkB
Xt2bmw8dlQ5lTf87fdHDzR+uVONKlSDhIy20YCtpjDZ+3sUR7F5iecty33fu/J6CO1QhqzWxfI0T
MwIwS9JoF1jZ44cB63L1QRYvpSX1In/xc+tMdPKBDZJDJSHWl5Swf5vZkgS7v65fn+V8t41e//y1
lz3k7ryKG1nou1tvxJ1UEbZ9v7CSp/FAJaWSc2eKsBJT0Ia9qlihTQd/dSIfU6dF9mz58+l+iV3u
Ivi8AIWPbSW0296ObwSVYtW0+Y7HhNPw9NC8YvJEEVRLfYjJJYJrZr2iEoSJ4q9BqJvXkhEdqg6a
kBMLY4BJmJWEFd+/l6PFnatQ9M9jj4QmPYhTWFyOnuPE4ehYPqMD9+wLLZxBVUisGzoykFlCriVN
TxmyIOrtuIRnGRF1q5uZMAY2ERLjfY1Kc0ouf714LEDzOMPPuteqvhSNCG4NxsnOajoLW8HOCWvv
59eTI8roRxbZy+fxaBBHp2kdqEbfFtL9b2wBp4XhBvmVgr8yyNVMVYS/vCk1bcOxqKoOyyaD3ZHN
YvxwnDLUAh457JrV1sju7BEOGJctLkja5IYFdXxn9FdJwRtYzxLylQN9VKhwZ8zx/udWYGernw00
mMofyOVX/ps6dqrHm8s9nxTT+kP1R4WWuUyUGcjHsWVXMaNdQBstM2+b4DWgDYGAxDYTHloBZFlm
mygwU9CP4vysl0W6SpEzKfzMfKvUjf1iw7Ing+TgpiSSZuypjJMTtp7yfFcXoK554bp1ssmRZLro
R60Y6mCeSX1aKrvOEmWqe2j0xX8VtVV0m2Pl4j2Cix3SmOMdmkVe+5zm48jefjXTrCSABIM+wMe0
c3PisH9Lu1H9p7JJtDw2VsR/rPlffUL4nFgpjaa+S1SYOhtAd5wegPP3KHHsFZo8fLb7WLPbvQLj
RYuO/3OWo3lrtzuM4Wdn87TFgOdZj7QvD6HHYBBi5GdEQooXjBDPetTkOzms2Panoi0yH1Erat5C
SQX8Hy1IR36y2zQ+UGdv+cFRJ1FWm793tInQYJ3JDrhDUiFhAYFfRvIJd9yroaug6vY8dLUO7MQp
NRTJod2VxQEBVQ0yoa6O05+kGYgPmnsXTGIxTujAMU1qgQrp0WINBJhFVtNIt1QDzVEiZIVqEEQT
hARN0Nf2n/X0rkzGy+arDsA1GGpIG/6CI3mQnqC68aU5mYTm5N+y4fWDY+pEUNAq5l3isQCovwMd
3vCn/2gfE5BlotLrukrwxY66ppH1gGGOnspX/Vh/U90b5scxnXptt3mNYEOY5shyU0CdvJYIkvFO
vyfYhYpJfYLqEJ9R8/XOLKKtpF4LBF6lB3uo+5YDO7aANRlLp1DRbzKcCG4g5MbjRtCCCPUcr34G
F3ra6MtO4FbT5xnLhHz693+6D2Srxa0a+VodguTHCGoVK2wsE5tsxJsvfWiTN1iq1NOGpqChC9zU
Y6wH3jsukHdJDl7h/iaNAjt5iHJh+eR8nYhcNQLKpIxsgZxFuXPwk3R0BBy3U3vKZKFp4+2VfLeo
d/43efrgBHtAy0VdzfSIrZmDInaJMhUPKDFQU9b5NEClS7eF2VV63FyCZ0dWz6S3F383fim4TRku
woBRlYXk7XjUSdOqf/CWca5aG92IE450yQ1eOsAWYWPBtyiDo1KD/FHO29ooImtIDgxCeGTufEdA
YL73mWcw0b+xag1rmH4t3oI0K3aYYyvTFcIgtoEnYnBgNgXeonFcrOCymVugJlPipgVwgXGPiE2f
FKJ0+j4hK5+MSbwkt2RTzFZ6P6TXtMhUyae/NeTWaoC1Rb/8wGydxtIIbAGZUfCex3YcXOE8oWo4
jRSMNnX1CBwxUqyCmYq7B+lRfFhnsHkkds73+oInsEdneiehZkiWvw/eX2I1L3XC8fnsSr1nO8eu
e6DRHOFt8y56N13f8aORZ9c2v5jz4K924MRWbSu3SbnalxjGZaU1luFZGNozkqGhGPojo7dbcw4A
81pcM6qBXdgu8SojMgSbBWdTjpp5VU2gdO2ld47dmmDBhKvIjBjnCO/qjkmlE8xo08gxSTXSWRAl
by1Nvwx9/EeCrcT2cXTL/hiWHh1UQ6qwoFhOs9WZaKjNsQmOaBv4PBipj4nDaeo4Lac8GSFTH3sA
7eMpnGeK1YtGPg2ph4Ss3b4kJBTA+iIFJhvaT4t7CWuni8cWi7v5mXDFvsm5OCmtm+erXDkg2HAG
Tarc+LNiBg9+JeUQCVf5VPpb9xqFN6ARWQw4VwgwITM1dWRpX8uhizJju/YBUNUYKaLf7SViL13n
0W/6m2PVMxQ103s5ubQ7fkSQ1OiIVp23vUHJ3/aYmbnABCu4zO8kV/vitdMicIzhQ+NN07ZcIctA
k6Ah31LGYZVsSakw8MybtQU2u26DS1uiXq6DojDaHAIVUMb5U5KYdj5i+yzmg9z19jkE/Nxxphun
S8orue3PckbzU+C8DUcQ5/4viTBs1HkP/CUfAzdBprrJ/1w1Nq+Llqyy6a7OBvbmx/KN62v8WiIG
jeibEcHIygyGmnmZmicSY/tvziuN5wvRCNeCqPQ7cMPVpNRGBkWg3aVRatj1HktjGI3IPDW0BmXC
4RJ8LKe7HEHry54p+aadOXyu8v4YAsp92R9/fOqL/rl06Nm9WqxOdLLPQzFldCC+RBOHnpdrE0h2
CCdSCsoG+qFy2fph2nBMNVUSfDIFLGO7EWJH0+AP7d3u0xHftfpEaLIUhpDB1dWVSIeX2eIECSet
zeKZcLBH0gOGAtUZYvCECsg+P3yynOWLj+Z2obaojpPhumttnh0nCRgyZpBVlZVI+BD0F5XPJnON
QTTvaMFdlx+GbGa2LSAxqtXdlEz0xccm74IVHjzlhMWIMhFi9R5et/pbMHdqG05NBK0B1nCojWto
QD5OBBDdMsApVNklx37CHDkZtGN2eE1FCkJhdigJSe8gIF1Dqg1n1qnep1Mv4zverfjf+DmVVvvI
R2m2Q+sQkw/8DcpWKeP/OTzhHSrZCufPRPQ0YnS6SEfl/QP+UOFD0gE5qpK8PmiWQCARy1/mRluv
3sfXOp1D6u5NH8yABCSqJUaf9mbPEo9al5vdHCoElyyMNgYNHtNlCZxYW+4pCCjy4+UUQ6c8Yai4
WWjmp9dH2Y8jP+afSqPYQo6LDnwyAe6/ncOb00L1+U1a3OuRnwk0SHIaVUKRDgSaToNz8WE+92bJ
XTn1z126CR2cMHFFXOgEqoGPy93xzxP3UFDh+3UdH2p75NeGsCnyIKDF+CCOIMkosnZnvQ0iZRqK
yKuYePfgkPmNE2twZbEAdYU+Q7bCRJ7QxWNQPyocefmm5FI0fSILtmPkvx5OCdjYaIxLxb3/1kTf
TQ1MCYWymqh7AS/3J6nzjqf6YSfjB2u+lW+dx2n2quJFCRNtkSqEbWROZZpCHvjL0elgFikUNXc5
M+8mdE2HOXVG2GIHrGqBy9fI1tZtxGADuTWnpFU/2OaLTHoCk0fmM9hrd62f2qpwiiTu7C//2oaq
LbEFKVNCTeWg5USzO+43FN2f46NhTJa4/2qrDRkFqnc20sD/YgsM722sgQytH0NTQKbcgEgZDHmJ
g72xAOkaoEJ4XV6e+BWLDyp68TJvUOb6XngKuxxs5rEFb2AIZiYkYOerQ5qMvH8vTicw3W2fcnjf
It9Jd09T0o+FzShhWHTZMNpyu75wE+N6djhx8OjRmO7rVZihSJFb759xlxeqXIqs9VVc6CIBHaSl
EI+u02IPsegxW640JCeI8FMrMHjBRnCfCc1oGPfZ+F0VBPDSWDTEytfmZbUtx5xoqIT74Cavb3ln
xreYQkOaZ9pWlBsYIEhdwUo321usHvcEhE+D3tiz32DOM+wcuspmvqjObj7dTwn63BMki/mNhp3j
ggDo53N11cXjx1dgey/7mstBgHwnHZkSdo3d3XkrUdNHZWoiFUk9HQw0hc/6XafuEVKq9uDUDI+c
V1kvGaMZCbzj7S1dVHB2m+/gnc9flixWgiwcR9pQm+vOVbfQqYpfUMoilukfe+v1tHkX3DnRZoW4
aJMxE0jojUbRTZGJQx3RwHXBdNEcpLzfCgYYJDvIf0GvfsXVCpH9T12RfyOcGkoDO8NFcXnvr5Ig
gHYqHRTVcKqcqenOfqqG7KRUeophPiwK1AGcg0F6li0NzOigHIBN/O4eYcP57XbCZNBRzkXhm9zJ
3fIujLgQnnPZqaAhdyizVAbkoAQrwT8ql0KbACt3m5LnXsB9MiBJ+IptWc5IsxUpznbmAvugN2Qf
ORp0pbQOSSGzJ0GVW83AD6oHWHkNGG+0PBGd9mhg72Qrrnbcp7UEWiEBGtyWUAD36ZNkHaJ6nZE3
l/SLv9Z8KnybQ2Cm7Q8FCTRtmd01gKxzrcs0+ig1IgC8bJJjdVye+WDr9Ymd6im0jse8iDvQNlJM
78UgrHc64FET9rqMuUNUG022Vw4fJR5Dk90EK1BZC4YrD8UY3vxGd35w/vIkcHDha09Y8/4+4ov+
zno2amNFglYFITDQ5YNxRHNdU9Vkq8zZVTRSneEQtCnz/KWhitIE/uYKsEl5QFvZ7FfpUhPSkgMr
hbLTqxknbliCfuCR44P9ft+IFQnif4X8ahlwXBi4+/kqkAcHhAVTRW7CMHnI8BN4x/yig3MqL4RF
zvHD4R/qZy8bH3/BePmx0CG7lSDMbA45VIJ2X4jM+cbCc9fAMPOWY9O1DhC1xpQdyBI8Ir49opyV
Ind05FLlNDBUqiQxqFrzpHYFRmtHspeAj6tDTgqu2VranpibqXpxwfmnpCsY8PdS1SQnLgkE1rap
9gCn4fuJJiz1SBrP86gg3kC/Ch116ccM27re7OAVGRnBLwV/4ccYxFZMWmfOBS/uLg4cT8qs7Deb
04cZW4SGJlbhR5OM7o5rksSB4d7Q/I2L3E17kBFkR0bK+gdqzkEPepk2ycVnmFSzuzWtcqbqR3jC
1zWb76myXOG9sJ9446UuCtP3LM9u3faRVdprYB/keo/dP7wjBJfLGfgOhin9u1dMIxJfqvxMsGRv
U9CdTrMjAci0/7j9d4t9gpJZ/5ivyyq0NR1M+5FdMYRlo5sGtuV9Q+uQqWgLYr22fjMunAPYDSpi
q0nZJ2VFB4ziseZr0XZUZy4C4Ps+GZFayHCzALhf1R5Y5JtMCOaIA2NTC1djHaYo3ZqPXd1mkQ32
Czcauszm5nASfq8i25u3sZbc19LZERJmFdW58yhUp9UByrzrWykkce93JELh0yKRTcKume8wjj4W
Wj6FTFAjnMHFcPrDL35KYWT5exUcC9yHjo07ATFQj97nBxGH7tUSsUv5szaYa+TtYyCnYou+yhkb
oAGV3i0ffsPt78/xRkxpn7cAclA+rWKYvGSaUfrEQssiSRqyKm5eb+QPhTDK2rp3752W43wqmmTp
dAEk1ashL7YBJDStV4UFE9hgWQ1CJwNp721iftYyCGKrrFrEX6tOQgc4VEtbPTz5DCZNB2JH1qnH
PrwZosN9FABbWrBxP8FBPMnj6c0LmQ0kmyg9mpOQ2OY65G4lbnhj/CQVqrvNdHVFzeRFcTOWMiC1
BCvRv7gIX5Fl4Pml61DwfZnW7vQ580TknEbSIvb1VECbfBgO1kA3L/XzWsBaY5HK5VjXpJzdMJgP
2oBaLivwOA+Wpq5qMyXosDOCACj36JkItLzAo83Ame8SW6wTHW4VBkWpL8IFBRogw8LXJtrPMOaF
V9cx/uHxmpx68A+Qjl/Fjz3dC7Jn488tfK87Iu8y5m16jrBSqBz/Ac/wNOW5BnFj1JAz0STrf1QC
sBjoxSkZ0FfNVbcrQVnwpX9F+IoCONPfw+mOSq/9lhzseLSrHl8sf+2LI7s+PNxbns/DjqJp21Si
Q7DY7y5aLzVSeJKe4dB3r6Am168e1rIirgeP0/btEbWIcwBAYhfpN9q7hc+/PzPYEHyiuoAP7LRz
Ka7TgwGFAYaPV3nQqzWHct104zHGcSrbK7cFoZrw5/8lrnR+jHxE9oXo/grRDrYR+xkjD+atvWrt
abS3PhXo5fPn3Q6ZPug7/3lujUKA+bxbD6dx8GbJFY+LROwl718O3kKz7J1nSUkO+G3YBith/4bE
HrwXPzNVu+DFggUwpNFBUrofugrp2FpT+hEV46XE2mUjbHBTievOpIDwckmLV9DimsM6xiVUEMU4
g9AxiA4IVBbv2kTB2WiMdBAPGnv2oodF+Bo/fF6nN0FiIWNvBrtqKLDrxKBt8RgwHNs0nB657uQo
XBbSos7sBf1wleA3g1J0IMvNTxKM6o7MDa/0b42bQeiUgDRlyHuFqIAj+ifXH+DXd6IpPrc09THB
IKFOcnq0LSxI8hHqS8csi26VReXPBpgwoLRx5ZXU16GAHoNr9iFfUDw6ll3VSw9kT6UTU+4xWhE/
p0yipV4ywOCMaTeYCGUrPx1LqVomwUbrujPjve9LARG/nuZwqTp2bZOgp9fFBITyh+QvCcWvNT/S
spGt6qpR3eJQMW70CfjqZ2MnjYqW5+va4yDiZwmFnITVpUxWc1k59Je+W57L1BQahvw8vWwhl7GA
9OmHHuEMJFXhCgKStpSAHwAvZCkiDBw1My+vrWtTXNGY1dw1KGsoL3amiH5pK3hJbBwYrgS/MJpq
uqg/elbS6oGNbJemdXfflZIink4Ejn/17esMh0UuYsfg0fbiaJK908IAb52i7QTCpu3Batxd7YUb
P6Uvk2fwzCWPBP2n6fh2CYpmxWArxAUGHi6vIEcGXJ+BzH/HEMPPL6avlf6A+HD9kmMa5Q2tSMJ7
krTZ0CxlgmuXhEaGkTY5c7yuY3PUvQG9mh1FUtcqMfVP1xdVwond3IJXhPKzEQ2pQklhGJ/dsfU6
U2HWoVODdP2zUEmsLk9HHPVovGouqhlz842yhQQpeS/hZkLPkFUdqfSRN1caFgg1Oaqdg/Q9XWxr
Iv3ej9FsqTxlKcaO26ULpQ11jAExZB3/sMro2RDW3TS3aPCU/SRJCR/hBuln5Oy8A1EAXBjfZNX1
0Muq5vSnWZcqvs7S5EX3z4ZhBXYPon/rhjl0xDS+pio2ijR+Nl5tBtLZS1h18BIi655WbBfOdCqG
Osttiz8i/wcnIS/E1FXq8hdlrXH/gtKy+ITo7iuzWlYqhpWVsDA9n0iqfAY7gpQ1dMyCyR08Um1m
n4rqCCmPJiPr5xrXMZQssgihGLOWIp9KsEiEtvgsn3HPsbqh2iIWowF1OcC3FK4ILenLekMl3r37
Bw/aGBuPElzruxdHaoGrV4YOrSWUwU3SQv6tjT3l9vGA7cOZIltAnmFZAS3/ZDG2cnOMOxHpRgKS
PuwXOpISIWcuCTo5xA3farW3NSStGe0nW1n5K2hwNnqoilcYtGC9Tx74hi0CUZEZPNU4JLeee0f9
A/jPqgyCi4Q1hCezXf0mZARIZNDBR+xwqlJjHTNM4t9lNhPo6f0DQIFZr0UYF3uMfGYuJgYMRbnb
yUyhLMxdn+eMs79bQqqBebaB1GWmuQiLFby4Xe53rAyslTwb0xL+mmhHU+yOREIPJfqEsk8eD49Z
6CbPkrJC3VuZoGWe09yOuCtODubYwLjp7/O9L9yl/F9xChuSxwSacSWBDhfqS8sWSbvX7H/N/Om3
LTz8pu6XMtyykEjHwCpySM+PIfNWP29GzLgwkoVgk3auv5tydBSonwr6Tr02mYOTH4NKDvYSzrt/
4hf0owRgYdaoMzqbgzyFdmJfHLkn4F1OgOElXkFFXA4OiB0e3T9Lwtq99q45KjDMSFQ3S01vKS85
jnagP3tXdi0IjbZpQbJIErdSaXud6yKpXdJefmYPCllq2P1joOuJUENoB0dC5abi1in6LsM002YY
q7t5siMCxkcpgLimK8ms086Hv1WWFxw9i8yipSB857W0owiNQMnkh/VOU7C3IWnitXSak/s3XKqL
VSoL72rVMJuawKtrPGzS01ygz4f0Jr/vc+NzbIHL2HUiWpX3k7Ri+cKVZSSjVoqBkQ+Y3a2SBfBo
CwDhUq3stp7DGbkn/ExA4D+jX9WGwxcrId2L8oZ+ycysG8MRVa3huNQnmq+GRZBJGbucPGWs2yVd
OGC2vUskmTzCm/7LzeqQidV2KcIBxbmVXsg44cqNhcnKOXsxZ3ynbGVjuQPB4OlVyraJpB7zNF2c
3i9xG7MTmLQjZbZKS1nVvvVZ4K+58DqKSsOGGbQTgYg7Fxjw4j+SIcNWS42q5KnkldSxCnNLF/Zt
HIhVYSOOiLyZNhT+T3yJ4INkyVvFvBp76XT3qausGxdAibFhU3lrPR5vu4pzmJVOlyUgu4cWsXyd
RvOMk66qPuJOd9TRnLwPalK33PgX+KqYVpWztkHUaUh8XjTVeo8NuEQq21u1WfpDYcNi6rmWWct+
D8RuIcOVal6sPZPU2qHPtYVlPDN8ORRJ+WWqzeiLMEga5A8ey2ouT8Mt+RHXjovQELmh1L6RZC4M
wMYvYXpwTSzkKLXE4iBnHM3s1GRS/41zucGxxZVm4KeWrL00N0e1PBinAbpMpZ2s/jd6h0OGfxJt
HjkYqqBGWH8EDIK9TKyDKmA2lSomjPQXW2b/0zhQKQK8WWrCHzhHg3wr4RIltTrdHPcqwpga1BB+
+Ih18sSP1ltV+QYUs8zVOHDdypcf9PUYVR1OOpQTg+JNpq5iYMAGfXzZpom5bEmhiTA7mecl2VK/
19yPMi+RvooYv+0L/X25m6YHCFT/9afVCfXVn+PQOc9+wA1qXoueH1KBTOYKqEedaYthcD9NxUNW
hkmS+7mDzvwi+eoikcAR7OLqioAepnp9CXuTKkaAcTQIqFNTCRKI8HGOQ4EOrGIx84U+LwitQiHF
j0n8GZwqWLJNgb//sg9YCpzW1nRqdMgGTbVmC6PyyFmXhD3BuVbl1SVktIliFvMa53D7Gq4Kvg2H
Yn5KRxod2I3NLDDXqrifpQq85SMi7OgoVBiJuhhKwRZnpG76Tu/J6wGS5p+Jcn7bSKV2ffw58HUH
gGlmpgulbzNa949bLfs34UFfNTDDq+EKYIM+d/98OfAjV88wWm0RYHDb9EC9th8uHRcSrrQNBKan
b187Rv2WBbXiFcJq5zYK4LxdIb0g2U91VS1bUU6tbHA/GfPFmQGLQQaCQlEi02BSI9yVlfe7vSIs
eENlDts/SWNwBnPoI0VlTlFdzTV0Bpj/1PUrrlmRRp3+5xGFigXKiMOMWyhkddywrEtrA5wwV9bE
As33OyzeYMzbCLyaSWfsQvI6PlI1uhi2FfYdb7KLB8tIaFx9H8FnZrzPmOPy+jFou+tUXImvFlVf
CfjyRIGVI4hZxR5x5jZVyPXHUNF3WPod5UzkQOyI0YMXh8u7VuiwLaMFKWjZSevuDyj4bCwlKFhg
JYEkcNVJlWLO/b3gl6ZgZqbK77ibXq5K6u2bHpsuYz8dtN9cAq5Tzvlnp+As/rxevFDtHNyuXZ1X
llQhNuX1Tl7v4w0Ustiv2MOb6RCGOAnBw67jtrNPTEpMmSUoOeNsPC6wUI4masapPSnqiobJ6PQs
ex/sZdyhyGwB71q1dW67/pss0+hjduIYTEy8cSkyU1WmSVrjEB2MSeQv4MuvzdQjct7IP2hKt5jY
BCQIlm/RR//bGRDIDEI3OMGzxP8rP3Bv4sJgWZ8jsaFHtRAHwf3WTZ7ueXGurCehrfKaTei5vWgt
hOQwxWxS5NhRbuxHE4N+bAdVraIh43nnGZp59b7KcGScq0BaUsIOl5zfxos8dbtzXGMTokdiNpPw
ua01WF+t6ake79KMlc71HhjGH4prQANy4YwQlGhuh+B5cC00T0bKujGA0FkzED3v1S/qXdpIn1X+
qOY9nForMWG2pP0/yLeMXnMgTjkE+0BKTXEhVRQ/VfEAhxcvegX721qnfqJxK3V6BhKG9mFryUnP
fk7RPkYN8uy0W21UyC3b2KjRKsId7akp3KwzUx6R41Lz2ykHs5KbktWPoHUiIrpFDpjzqWb8AjUb
7dM2O+LXUaIebFts6KJik8sNL31GbdTd6baKYAqaLUBhPOAUyq9O7R1s/nzgQmbUXjyx+nV6YTTt
+GYNBHaOpV2yt2kJ1+c/kbQbI72tljV88Y+WoWd+xyjHFmQRRCNHL4WoLk++70uKMVu29IMzs7lE
Gp0XYSsQ+ofU+6hEHlxHr9ivErxnawJV9btdPBomqgDuqu3dORF6tCgGlZMYtmf10/U2lVrmqiVP
i/UMZDo5GKEf7+9SbIxLW+nUbFmogYtfr0LwlSmGoOqnZ1rzdf17D1zS9XqCjl9cNAXtv92nys8A
MtRak8j6PdPzTZiwxyqNW4SO7rasEzQQvxfG9Ji87xc60L7goyzgR22ySaBR0ej9cIR50eOolJcd
czEInoU+cWvmb3SHXt3qxHmwRKAw0iz+XCElQruOSeaXKyDwwcPaIi4cJ15GjTuMFrI7sCyFIaZt
Xr5hE9ZaX1ffUyYZ/He6EQDJ2jzYtV451SRfIJWRkasrzHhGDCAnh8FyPux2meJb+oTdTLxvgHWQ
GKt9Spi43aG3f5PZWRU50+tAShs7Eb55U1v/9mIrrUYAAS6/hiJ+CY4JVn+fwBAeatjveXmx/ekt
1ltnmncxLk860tYVrXHXgGt1CnHBahnKC7i9Boexv/2aX+kagi8PeC2I2iLGiKnx2QxCVMMRGkcr
BovkKjimcaUOTcpd4Ao5sGb8cVparHpEiazWxs2dbbJYv06m6GNbIUeAFAOtETp/zuDRIeCOksdt
NwduUriNtnC78S1V81Rvc2jiV6PyteDK6zdmYgljy8C9JqDgl3l56l0RrT5fEx9N+LZikS8sK1f5
vJfhRkgRKB6NtKmfNPWRGmBbgxbrg3LdwvF701q/EmVe1KxepuPBJGct+u3DPoWlU1d+3jrn5c05
1fub0jTHS9x2CYr+Z8KGFsAuWYK9c8q70YA/7bhgzaa4jmvnWz/e8n/3E+3+9uthTb6WZKUsOapU
mgJ442nZDcKGLsbMhrbj57jlG3N18nv1Drk4Xiogl+YB7Wks7dNCOZMAZr7Gjb3MlRIDqp4jaTZT
i++sAN0H9N8tk9bm05ej/CEfgLvxXCio8+8rUnNJ3BplbfolSJYvFgM8Ygv+mh1D/xvFF3fgfyBD
RPgy3fOC/h58lsecQt9KBWzk0d4+EpC2ewuCrojn/tFkUQ11sbSspOc2d3hbVs0cnJJ/w1KIYPtd
OIsWliiJw0rYPzx5ccH4QJ1EqB5CArJOqE9w6k3hCEImimeV60zAFIfFIlAKM2a+YBgs+OeRtPUh
z0xQAOQjQvqROu4/kbsMj3yETOqCrTL6GRS6BW/VvOywITpFjyOYlv/J0/iE7FJloDNCmTmNLy4X
wPkwcmQkA99mFxGQ0kF4iQNWarct1690xqxK5gfKg6hxxQOn14H8pvmf8aIGeGN/RKApjd2nk8HW
lYDEBIKBOXJqZJF3fvDyGPahNnQEuF2EG/COTfY8tclwBTwqqPRF+mVUgiv8hNujhcs7bNGpJM94
+vu+FA0G22+rWtmPRoJfZF53mJJcDSazsKz3y4KLesL99v6zOg3xwqvKYdCdnODnvYOdj+3JXyZC
TzrH89M+k7P6CILZva+M/3HOjYRfARKlrsPceu02MMLnGmZRXBQrAXbj4Dmnp04F8kjGaHTNyatU
jnIjMkteLr/3EjiLs/lSFomoDrqlYVInXUKhaaB7vA6Opq45JtPg3WKbH7v/wjWbXc/FSmEFgw7k
rTNoSfAjL+TDpvQT48iYVQHbK0Dac8KGUL6yKoY39KztdQRFHECqf8RljMdqTHYEHHxP83uCiLmH
KfO5JFGIyiewDB7Wdm3TThEkBZc4l6c3nJT1APS0XAUaIL/u9I+xkbvXW2AZwHpjtFyp+0r6hq2H
OSUuoMyDOC+th1iLoIRzjUcW08NfzmN0iwLrTeDo4Zfa+ylgZUancjJens+8cY2PM+oYuPt2MPtK
26f+WFFmzLQFufbrix1FnTL8xtXTdSTo7qwNgarqtT125jBjDl4b5DHpE6dIiqiXwKkHAZdI78Q1
2+DZUr+kpo47FH8F1ac+vAoph01ULYczNFYQAidcyr4B9zhu1fPhcMOtnxf5wUEGUVPT6SuQMiBf
JUBEq7mnbgaQaykYeEWpihxsvE0HBf3iU8aw/eU6cSS6wak19At9wdPGOiLNdHo+FZAzF3PPG200
KQhcBdG2fKZisTtWb61hqHuMTW4XxjhHi0iji5RqlktDRqasB8jeM836OrKiB64V6en9Qiw/QTH1
6a30bPF8XaW0rfEB6bMbTJuY/azBZ3DXXDtRmzlPjiKshH80BbBEdvvkFwYPN1rqKNH+QwSgsAGC
3wGbslN9U1qG6j1MEm1MgiKCZCV6EKwyYPFhSxJlz4048pdSYl+HFse0Y7O1HjbwbMS51TnX9M1u
rP8qvbFO3CTpwHhf4LiFq7EpUZM4ptbVh2p2AIM8xJeu0nbkS9SxKQaZce2LnPA+PD4KhYm8PNiB
Qa0bl1Rpsp0EwG3HfEqKw5JPvYiJ70WvsgwZ26HyhlVG0+HoCm/Z3kzVqCYllWZct73CH5RJznU/
CNp+Bq6/vF8Ry+xR2DQhzdVD3GHsvBxrE5XC6iMhXJLJTR6BIEuAMOVGYiS+7N/6m/QIfBOOfrhW
5dL9jH6KlwPdMAlTIQajlT6sM+8TqmNaOIJgRmt2i0zbcZ5WpQiZi71VgsBdLt1qI8aWZBy3apSW
O86ZIE5TWaMxGBb019jSDV//3WWHgxXBMGlFbn06CvHflmBCh1vtCLPj6GF7zT2gbKD/vl+VXm76
xUgPhq+V3vqvBtP5rePQayjmyeigFGHk3AWraH2p5cSs+FjyHt6dGFUHtwPCuhJOTVywu24sxiWR
06RxpVFiT6O5XM+kNA9gxJVNHVhhpKZIKA9wD44Dok0+w3+7KeSVay7cd0/xIRZV9+i6WAxKR5ED
iZhzOX41Ea/0PL0C3ZC9nLJQNtYPIfSFgY3EKK+XwGxmNMJB1mtNPtkQ82wqTgJJi5uuNrVCWhcs
qsnWMpOmo70ywPkdKI+OR/idnEHbszYIIaw9Wb1gLV5wuA/DymJReI67JbOm1n5tPZM0Kb7s8Twj
yB75l72xFgz9W7sV70wG6lVe7OgC4SFJcjB1CmBeRlmLszNgyQ4bab+yKxqIBXHmkibv8w54WCZO
T6PWssNeikmZEpbVKKGSSfE0ht+rIO8W93PDpQqg9vzDngY1vAbbNkO8ldnz+27Qh041MDGsASPt
Vizt3vjRsUbqEWeFLaE8pRm6HYDj37OWbu6rnHiJqOheM9qgBYqoiRFljv5yIGGuEV9f6VFSGd5Y
luBn2PvzR5/OjgfKTs6ELY3AFZjV1UyeqGx39Ny/eVMmlB/251uBNR87Umtv+lThQ73GwZ+Iypei
lbSRgIIzdMlrPtvwHawoO3apoFdOyZ+3qUyhqP8SlOhldcqNS4uy2oRQ050S8zEVjmvkKt3Q3upQ
kYvk6tExEq4ASJWAkEoTgF2+0rVHfr3i/qqkklPpwTYQ6vzMLm3R22bYWYERWow0NqqlrGkXhJB9
gAfbvoFRfIS1x/RaV9xSw0JIFpLPnzNRW1SCKMm7jhPQZ6WHH+FEzAfB++DrJq7M/JTWaO4+dEbB
GGSyq0QjHO95MERehC82t357cyx9BzP+4LB5s8S/ffHvZwzLYv+leAaMs+91fajxpvzCfsvnj59X
R/qtGh9B89subIdxtDklCR18Y3HwT31Klfru/T9vlzgZ4Tt/pQpUjd4R3FwNkEHljcZ2m8iBgLtr
SfDujc4pFb8jHnqOANkVkDp2T2OSPNe0zt3mFHktOgj/hes0fwH12xVdodPGXjkP4R3fkAcY2TXi
Xwi8FrPrJ1mBapcAxmqR2q1HtLTo4BQf4v7g6jOTKDERgu1aFsKfTRiiNyjhqQ0Ge49MwEZA4JiU
8+MNjm2WphH8ggcomsFh9/c/0/ga1E9Anhqi8zgOUPwbwSogwGzgXQxF74RxU4OJiJPqVRD1YspF
5dF24Z61J15EpD4VXrtpf+WejnAWxtnlLVwfO0iBnH1nafb6luNvDsQK8AkVToQURCORtmyD5F+D
YCDyKogrdfh5J/u37tlhe9qqwobiEkOBlgDe2V11M+scg0HCqcDPEKNbynQHI4JQ7mtqdoQxu7Gz
PWzjUJQilAWVgYwUdeUMB6cT632sWvD6/z42/A/D9GvZ5mjQ31GuPo4GVxTr4NFlxueLkvAC/0ds
a14Bfsh7ePJp8hAosDglvXCxqyoM3MkxJLYtjxmLLZUoAIVxu9TiMO6WPi4tsillmENhbaudiDB1
6ahg4lBo6Y0JBI6d+hutCR/66YLVtpc/kdW6+wf4XfImgaPoJEuQgrzN5JBZT1pqrQcxNaHewf+/
ZlEdsAhc8sf6ZPwjc0z6E3oM9iRScgqG88trXqVt9lzl6OHgZN3LDRGdvrrSi543D8LdCZjBusfx
6T7i50oAVtWeXNT5AfU5UHzv9zHq73XuKXDuLL815lbNyAi/Zbxh2oBXggD/738rHstUQfWCymxv
42+b1NGJKeTOGt247ktKV7UadJkPOPtcBXKagFPhtQ+QmQupFfg7ZGNAtm7w06zlRTRk3ZufHOj9
hc2hOaaVW/hREMG6h3mGjdr6iiMZ01LqsEGBEzKndwH31NCbTFT3IWXqGyySVgHI8a3u4WbOw8mM
NdyXql2QfeLFFeJ5EkO7kQivzA14WNRpq/0UXAgGKPvFUt1DlHqLskVtbL7PektTTq1eayr4wx0d
PP2PBwR1sdhefvLvN2YF9RODPMwLNIcsatacLQenAxy+lw1Z6dFFf8mdlU4rv+6jll4XzGUrBqvY
U0mf1uA4jhgl0V0rZV2cXq4ZnRUkIrDavJNpw8n6vJDuSs1wYwIqb0AON3pTjFlj5rZ7u2BVVOOd
a95LXASK7P74rygqZ1Es00JhJspCBX9AwY7ujDtD6eUAqr+OoY9ji6lcSTgCblZ+0734knzvBJ/u
mISJH1IKiupqhlzHhzn/hJ41X442z3aJr4SAMq1+xBqiJeiy/PI0HeNQpXq8PZZJlxItl9p5jyu3
/3F4/NyrP+xHTIh19irwgaznt1mXcV+lx4IpuBZw0MRjYlt25QLiO4o5WXU1avvIK7iZdU44hES6
lJMNLt5MUD6QQzD+6zRpSoJbHJr38t/8rswxE0LGiP73H0T2If2FU3Ha3Gk/GAgM41pZI7l72pBv
pO0w5weFp6hmwOjsKMjnoKkf8aCN7Xjjbn/j1cWCVsm4H1B5at2v1FrQpP+m5IkAviDtnK5r/P1n
v/qUCyRkCLWG5epGkyX34bKwSxqEvCjEGMSjGnbjCjukOE9Y5jhAxwW/SuH4f4UCbyFtVhFuUF+u
6rLiW9F6HNcpfzmsQqMH8jkWUgV8+AIpIG3qK7EI6w+HGxdNd1hdNrtNmfFNpOkyW056xS9Q9wpT
3H19pEpz/br/fpI8PxJYGCHe+eTJcBSjilOJ3Jn9BkSHzAyCFBV6mcZooqi0Tn6fJejSQ/XLT2SO
wt5KOOxX03M59yvpZoEiViTOhzHfMkmRN9ZD1b3+nSnadcuIIwlQx58IEz4tBKYwVxM7N+1qA8ef
V/HXVuryDC8RWExlLGiRGw0bC8zrqoAderEdL5ZXyDc7THGzUkpv8zKVOErXTMUIkC59ILNFy12x
EHxI/VtiHRPelH3Hsa8qZVKe6UDiGtD4q8Mqwy0ROJ4zN+cFTb9x3C2Nzg+CpJOrPbuUjQnzXPGd
xywLtFHR9PJb6YpllIoVKKSxDx+8MfDggr691HnIMsyCANYKx80hKh6u6FfIGw111iqoVSh39D15
b9G7J6OXTOBpdXjzx0mO7j99O654CPYBIAztxx2CoioPt23mu+H5VKVEjuezkbTIGae300vnDYYk
FJhIGLMHA9cTOq7MSqS8TZ83z9kBOcnMs0XRbAu6UbMrkGs72cfCb2/fIdF+CHVwFzp41i7aY7Fb
aOZ3M5DgVi5RpSG8Kz8o5qHfDJ15ojNL2hlLp9ZWtIEtgd+vCaOm5gDB4I4S76SCH8nqLakNfC1D
mWljnbjIN4aT0fVzLXGMqYjta63CRmkw62laekeDu31rmlhmPvCNazCkTejzz0rGHBj0PiFyrH/+
TVPHlPTLIvWXzyCFPuZd5eRMg/zlhYiDFX+r6WsX0BCA0uwC4TygEdHJNy8FPOBOpQ2NfUPpUjxk
SoiDHf9maVaQTBHbO/L96Lz9aIgXxutlL1sD6qvjuvd6JxIt56J57ghqNL+q9EmCU6mJ1/ZBS8FT
3P4J2vcs361AnuEK/YUHu2rQg9eeoituNq+ZU81tXBiNE/Dqm9xXr+mSzT6e7ieoJSWKjnyJzshA
mJe2g+8EFanb7YdadYMbXlPSDN2OeELSuYoyiQWVc143cCvGk5Xz2N4c1dg/mREb0yUzBTvHgzpL
fvlvENxvA3ObpA1RQbFSvOasQvBT+mdWOB6NQoa6zgma/CghPoa/wccckReaDiDqK0mPVHSrG+PF
dg9SRx5+yx38eTJA/CmcSHi36otxA9+dmuo1THUQSkcqICBVzso4jTQzBZdIs1eHEUW//F41BG2U
DRGHIFX/mGIkJEXbyxPzlZ2B4uKeS1CuaPeHHtKkVwOMzHUlI6VNvT3xg+rM6mHHZx6PFMRwaKQ8
wycGa7Z4Yt7p0EZ+VsV80xhUej3Qu7VmZzWP3k1bjyIu62E1PDojCOrc00WytVp+jgh/kHukJpYv
4QGkEUej/veFhqYrUpTO4VarPfwhzSaerdF0rN9tnQGPm4QuFF/DrzYCvxKd0D8d/l459C+GoY8m
0d8csvR7aUA8DR7fXVwBDRnxI0JLIYEYd1nGAdCe1YkSiJDzqT9jbjS5ZC13M0Rsp5b/tG+H8EwC
hZNpFYZ/hkUVlH5/XmmEox7i4gv8nir7TAgFtY1Q0bZCaxCR6caywYXdWoNQXGVZqk+9LcU557hy
CPoyP73y3vQoqs2J6xbNDyd/i6d7dMbge1TxveLn1/Y15SeVNiPPa2nbdfTxDf/jCtmeM1u+bHAg
JG0JZvK8iOTCeQQ2OiCBZFKB8RT6vpZiIYhN+JcOMnXNVcH6a58DydmPnDAvEHmkkVx4py4s0Xw2
u7YFK1/8XH5EfzQ4n/dRu3IU+zXzY1OEgxyB+j/ckOgAz5L7r3QhoBkqmW/GBVOtlFrh0N8NyaV0
UYGPtmS72NizQCVd8R5c3nE2vdfp4QJViX0GudM4kM6IEQYA2D68JhM8iJWgiqx8S1OxIK0I0fJp
GhW12CmSm5J4SwEwN+dIUn49eV6UGejOh+EzjrD0DgMQUE13st1FpuvTBEQWGqwDJsyPwHTEU31L
IVyefwm2ub7BzUmXtzVd5cIBSr5bxa7b2UnwkytuFuBKjqRFRlfiwWRkPi+1H3TxA1KDZr7Tx+nP
Dq0tL8+hlA/eCQEjIQU+zAk0RanTT0EamV0FrJCyRrWJQeKNXefCBziGzTFi4I/z3ge1WqpfnvBT
VJ0bzx0WI7W3kiKfZ5MAfSZUkRYCTuwXu+bczds9rEf25zYuqa6Rz//P7lTztmRnDp94sXW2YtaQ
J8uhTseEStSpi7JzVV9R9UkAAs5Gi5n+3Tm8yAoVRsggRwJYsMRDSX9KWhoRcbYhDpy9htpRPlku
8n7CW+KhV7McXHX68Y10MbVMXp2JpcZxeuvxqXX6AQ9Ni6avB25x7Gos6J5hitdMFRtyAVbrlJt8
Ywgqa5EWAycIXiFn7+oHGoXHu/cLnEZQtdSFlF8wP1Xw5/KrfzdK8l5OSsxwgkm3WnFBDrHYBjb/
6ufhiSQ4Y3mBPVt6DHGrCO0YNTdBAtrzjQW/8sjoUIENYOGTNdqzGsDFU5ZM4T7DDrFq4LXUjdAV
F7rLRpqQgGm/BiDSpJDBypfsD+cZ9OKu/w1OLXvPvEWpQFD6E4qib0XUohB/oT0aThiy2Jnwv8hU
Zpd1ywoX+kHixO1SPeTcW3QbbTxT6kxUWR1f4rNUUqIWrzHBOfmb8dlMg5b5HxhVQU6u8Pr05cAb
4rrLBgNTShAPtsMhpH1RDHr5+O+v6dfeX6nLUoxza0Idx6VLiMvTgn10oCTxzQiwMzvxQrPvB/T1
zC1wz/LZSfUcjP61kHeBApZ9gwKh9M7u4oxuONhHM+nBYSpCQVs1Ph8sr7fZvDAtPBVmGV/WFpV2
0xVbsK0vXXe7OHwxWg8+43HLmUepFJSTnm1KhLwHgVhjg+vP9hANPbLe5d9PFXlfg+QfL1v9g/nS
5OyQg1j205pTU7Y0GcV4eZzmAFL4rUxbwl+il+OyV+Z3hgQFl8t2JtjADPb1CfY5onKbTX9sUjk4
27FFiAMUp2f5JWTVDUuU6BViWaoRdGWrLeHVnChcty3fc//7H8Oj31qO1WdFM5S3K3+YwVZAXlfG
pqUGG+YiJnQdzN3H6dHmCi+/ZwmmBHuNYT9RDzBM+Gd1O/Q3o6qHOXf9aibHFE7bSkvSbC/r4h41
aVf7FL5lVtPrUh3NTtiUmUqPfPnptHUB90FJOENZDZSTrsvLqgfSsxjod33DHM+Etgrbbf6WEox2
ZFpzi+gkCk9O8tqMaERbJVrRK5ZmmN8Ku9cKfMHZ2ZMM/uot0xSVwKjIVTtO6fiQ7ip9jYv4vRIq
34pAGQfP6X+3gkQEkRrmbJDPmgmcO8p0GSMsxUtEnN2aBroFWoVz5yvCG8OynU3eVw4TLVJZZ17v
KPLxsaxyz2g7tr20ircYZo0MiJNzplqSm1AKKt0B+Ccf0x8pXrGDlsPaHl9DeDXYDwSUhAEHoYfk
bKzu6kBohF1dnLaTU90jLvk8zOvtjofnXlS2Fk2RYpQ30eEpF95K/iU1Fv+zyjJZNdXcSCGbSEkb
ZzlMIHFLo1Ie2BquPpU3gZL0doVeR6qyvGMr+P5y+kk5Md+2a6G+x8LhTvFegl9nD+Ln2xfSEF0E
EiJfYlhu7i9d/XF7t060V489eBm9qomC2za9VX08DDfxrYEFtmkJdQ5lEzA3KhiiP88SYkKaV3bw
vf8jf8SbaL0TcEXbukY7nVWvfUkuRVTvau/W1UnRn3Ub8eoRooUNJCW68BD+9jttIfzT33hNNv4R
w07qPkLeKiNUpa5+F7go0etL/3MZj/+EoysNTySJymyzooHilB2l10GXA/FMJtw8lc62oXcJtHf0
Id3ntRP52tfefEZhjWtdv10ByZ78u2/R9CaDHem1LINr4mq8C9uNSfmX92PvUgFdUJRQd7WO5itx
nutufwQVMJDbQNMYxHwghp/SoFRRtYEVWE8Q5Xo2EMt+Ek3wRrPlV/vsdtokgZnrJ/IoMTsi+BoN
/4Ifjunb0OKUJaCLycHcHy5J4PqDFSoHYzUXF05cW//ufN94N3WNcErUfEfwObFe5dspVIrBiX5b
W9sQEV57st0/VSHsrzsIbWNVHptWN/BXENjmWgKF+ZuCmWsmze1Mjo2VRK2iMvxiTcxAuJm6lPoO
6/68bLumRWr/y2RgTJYKzE3XGCdEww8SoHRU76M4lWZSUCkszmu/IRi8y5+DUWudcOmVyELWjkPa
1UZHaXdcFJFf15xqZBFbIhH1Wm54rhUCB8BQyOYP6VY8h7sa5OijljkLZHj4jVvi82eNMmuRKFgf
PhUHLrGyMQ7fTuKkEPfrH2H/kBKJtN/XyvUDqhIam8Zj97GDrieyO7/QPUcxcdZU0TyIuBbt6J1y
FyfLD2DT4pxjoDU9Rn49jDc2omWqHZhgq6o9I2ONjukXkYjSp6fUjWtWYf+ZsEYWxkfRt/dNbUGx
J5wY9/XC7NUzmmCvHF2keUrgdJz9gU8h07cxRoMZX+S+zQz22MvnSCDLCCS1hBnDawXbV+LtvW7R
YEZtj1Yyi3/ajjDNZBzm5z2k+wjiP3+EVBUV+BMhCj3/Dq0cLDQRTyky/hfaSvolR7rvntYGT6ZY
ceSuWVYtA27/+GeQn4lGmEz2GR4xlti6x80QmKjJ3BSX6Hc42zNzM0Mi1ox+SVx0WWKeJxawLlhK
rmTIhx1S5WUW7GaitD5cOpjQqFPqqIwnXhqzKtt6RJomj2B7bl1KANERjQ2txfat7BZf1NhbXzds
oqb0Ew3EKxTkK2hVCJOrLrxUlI8AuCcgstBzK3TN7PBROKeqYk6Co4bUkDpVZrbZ4IGlGQMXC4+u
D+bXTdx600qVHjkYj0ilmX4ANEQEo8IJZkGg4e/anQ20aL7hLqLi1HOeIOwdI5sGUIhdd2+1rs+R
Do79NR5b3e5+uNlhkgjRdu0lTkxPprsWnCMjcgXpr59XKlWtrx4gnTdl+Ly3VZNGiHGfHlJihHeF
ygS4Jw0SCxDAywtL4gksiCLIw1EH4NJomidHcOLAihbvI2/M4bb/Ml9J3bwrBGxpDJLWqyg55h/5
Il0NbSZAD92vDL1S812POXM1a9AJN+jxEnDNZb62IgPh8ObxhTFp5D5rmDjfldstwsc14u6BMpoh
sr0bqtJVD38iIDE7VfxfazPQyj4skxqj4xgPaOEP85ozQzixggtPn21G0K/EPHYKHXqyYOSHD6cd
lNYgzJSQimn73p1VJ8TgUgCWDoC5nWMJy31Izy3B5YqZ0tcEHLY6GSiq7f43GjXBaGznqZg4l7ez
HXZkeiSYp+DuNSZ3pyGvr5yMG+VSkT61Tys9yu1P1HVngq3gZrwy1nGw+RQoeg1qhN1KOgIJUnBw
bOY+mROnDcBDDvSXh+nB3Qr5dauKcshpXDG1Crvf8Cu5CoNyWThMJYqt0p30ds7APoDlR/3+ZcNh
+D4sfSmgZOZ1rkMS2qKomrygKPxRRT5PSU6Tid93UiJhKQnQY9FfPycHIW7hWrxDW38gy+xrKrZd
ArBfxJXRHbTBO7xFakntv/WaxrgBpnbCxE6SJ76rpgVWr0k2VkDiV69sBk50ssWTT/NEhqckFiOq
3oRqIKEwyjyrl8ZitY9JNd+DpTE4nO5ur0hW5TjyafQqvaFeFQsNOQjplYKzdO+VbynHFkaI8h+3
aXy10ip2KqQylvR6lGaCKL4N4fJJR5iwiWUcPuciSv2WziknJ+g5g5buXDLfL65oexokfRpexHgw
m5I/fAsQ6L0JeQB4dxmDx5E8wbctoiumfDHIDga1RoPKAN1ZQSb2yaejOwtKbyJnV0tDBK6akMVR
f3hc61BZtyFvPMK8J7CE6xIsa9/D6muGklfqMMrzv64phb/KYoRxR5SomnLXwmeSD4k8+FhLZXdl
285nCmTPjQdR7FpN2uZ4f2NHaevs0cID2DMNlrJk1DvHZvPpaZ3wJsmMspBu9eWvFhdY2VMHfzc6
+qvmwikcbDAJsjvm6EaQtRHOv7XA8Za0DI1hB80j+De4ZaEOBJrJdUYTOBd5NSJAdajA/iZAOu+F
cqQw08bJYIA5Sj5bAOpiZtNYVbpzEv+dQthYVJ3sY0U8rt35BVnlV4J5mytJyi6ayV0iKKZ8nscb
Ynd0gKOg1BkK4YKoUI6V6y7nDT9LBvb0FYMM3iuE/yJGfpn8PBk1GJuc4v+Ux7t//BehnzJtGd0s
Rq9jCCEhj9AXI0RvMEyEw8YnJgfDiciqQkjQ9P4qW8XR+kBIGhWe8Goi/k/RRQ2w+Vn8YyAUi/pi
7hZsMRh4eURMG53JOz8LbRJmDgOS5oRff5x2pOplp5abRTixqIJo+HPfUx6F/iWRatixcKOCjz03
K5/QTx8iwcxWuTNvM24PXRfEUVfulttF4x2A94uhtfDs2Cka3luxgTIv9hivzRck/O+ERAuuVvYR
buwuQhbP6ldcUBzZzuugd52soD+00P4PjJZ5nTI9hEqrW2L3YBVKNjsRND0GGUWeW8o0xreLO08u
pYKon0cjxuKAVlCm4F9ULxaio+9XMeDrHgdGBkpDh+fkJO15F+Y363ja/HpuxW1VtEsLTPHUjOqm
G1+gSR1M4Q0DAX7KjvxZH0ECAJw1pi4BPRogUBe9F9SGXWjMuQrgcjK5ONSfhIr++/4Z+ehY4KpM
UTuLOMuzCl6vvjpnbQE15PjxkqR0R1Yammd7cjUswpGLOIXzp/f6NQuMcQWekMEOsqMcbhDnoI9C
OemJ7UbB962dvIBZqo+eGyTqMJmz+sv/becGzwmaWhtAY0ojKhAPbqwY7P07IycfxTpPmqEBtAt/
vLlgNfYXdBeGGuY+mjD+CLeUQk88s9IMUERptRWm5cte+aLApiKAGlTLvkm8yWs97co22rkGfxvp
f4sNxKVzJqwYP8sJu44mrtu0M0wyrZWkh4gLV8ocRgsaNPxoT6E558uM+rnecDM804iRwxuSBQfh
/BIaT97YCXQfoPHGVrj96GoffuHfMxeNwIKEPssOqEFlPvCPehPC4R8zd2TjUtNb1xuuT8fYPJhL
c6Rxj3LFKjlCPHMd9wobxNNiXCs1xLbs6EQLfsZiJURhkCoFL7RQvIqXgJIGHrF5J8LFKtguJX2E
9hrKJ0V7t8K2YrRKkMHcCcoXaAKGmT5ucqfa70pR6C38OClpI/BjvLIj8YgRvcQBr2mP9O7aS/Lf
vZXF3jvYpsuCjSZNmUrDzDXxsNE90oDvwBRJ1crpzO2P3YjuYIxk6LZriEEMhSb3RBe1kQqVYOsR
w6U2XFckPnUDsHAg3+Mavyy3NLAmv+hDfJ9gyYXfDWL9W+Z4cgBOZlJ7c8xeLR7QAAqF6TxlFEnB
BO1S/z1MCQpmfriUY+fEIWu8mPct05X3KnUIJRDE3hif1ykp++tEedPXauHZi62+0v1SnbrBbuFy
0qrk/C0W42ywgbAm0pqWdwcb4uBkOnaqVGbW3WBPod50Fd8f4V+K7WieFeDjfx68v5ECBXm0jY4n
PTNdTR/2N6q0ZOv15JrYyhxrlzHSFNgjE6iOgpvHu4WmvL0RyD5JFXgnYdfziOfCKYXTMrlmuXsf
wGgX4VcOkWRnnPIa4gO7ex2eF5QQgzY8q8UeaweNZRtGPeI19D7CbxhSJaawRlaczq2KN9p9zj2a
rzs7nOZJifx0E1cIeJBBAyXNWTSN1w6ThDd0yLti8v2BP4eXDJUR9pZV9B9YLWH2VAHKkIQoFesk
Ozz+VDtZnoHdZzybG+6O8NUyS9yNnmIlCAXQbOomSu9aoH5rzeKErfL2VGX9V1w9Le/mHCqzV2Qc
HaMUKB04ztfhfwOwsdzoN55mu/23bDpiXjn5S+se90vi4ZRdkdCmSxVnX/Gi01Z7fyQ9XxO0/aWS
W2hTAiiWnm87EEUeDBlvKDIbRypO87qsndT14GnwgubvlK4fGNSZ4JPLj5/MsxQ8aXquoSxmXLYv
uABySVye5gt4Xjxbwb+zr6H4A0wpsBCbgAfTJ7mOP+t8Ync7KPwYtwcuQhT8I6dMh9qPo8su8aaA
z8LeBofaCCXFXW922rxaX9JOzhBNHR62zNumEFrQBTjtPOrcZ2mM4x3ukw7jbbdYF5vbfNsxn+XR
sRozOmNq0/Rq+zTNYFBJ++wLsMvZ7TMRK+ToYBfbN1uhxDMP/TIHESD6L48XjM7wdrwURd42H9w8
58hRFtbR5DDd9encgM0Hp39pIf/rtYavMLiB2IaJ6Ps2+XQlhCyFXTI55DWMyLvhmLY6wcI5UfEP
DFbNdJNjJ6YzVal77vXsT2RE85lQsVYlFSa9X5vYQwWIgleLB5IS5OpCf0FMa6s9V0Rqi8u5t08l
eVDgNbshGW0H1VQPzIubS5AZz3w6OTkHYElThHgdCDirwmcXGsQLEqKmYdeIhEHrKAuleGLmchPQ
0cRyX54BC65DbW6C7Wb2qxhbDCf1oncY0pohx4pjbkt9+iFHUnwvMbY9DLVPdvDBzsOmygR8y7Ox
ag5b7Z8BhlC00QjcvGx+9fMIk7nszcit+c5zXgvdiS/po1kA7rk0cgFsAD8dmcsUtUYu0m1+/mop
nbUvav6oaT58Ix/hiSlRxHpQVFPe3ejP4uuOe460lQAZ+1t1gLbYRm20W4j/ewaD1YUcZkMrRoQG
0zwE/kw3h7LpiKfBWtI/jq+d0Ppdw3MdX7QV9swgWPXNcmgAZEGd9wNOzTnjX4zjsZvM1K+ZpzkP
iV7ez62w6ErfFL1c93rB1JQFXc6bvZmuLY2IVJ1+qVcPteVxhMlzWvprLqAq20qeeKD7oYdKQ+Fl
8UQ/iPf6ixwJuPSCskCPXXvDkaDcMmGk9UtBURfifmjOpbPKie2Akud43gr6OpllNjed9JKsYi/H
fS00YGFJhSMLP7/gv2Xlap6HQUDrqc8DUHUO9dspKNC/UxCy0b+bI3MLm0orkMpviWYRQmfqZNUu
QibX1nNODjLEFbQ8km9xvqx7G+N6pY3i8TvchmwMEYCG0K0UngPOnbWdSxJAjlRluiYvUyQklXgC
3XlTDEYFxFbmYXXtGvyGxQ0be3O+oThn++5hvIyGuiRiRTo+IJz1e9gAjhU12mQGv2Chqx1Feb0g
VpRzSnEXQN5PDijDr0QsRqWJAk7z6rnoSwDsMJp9bgV/bgJiF5WRUQ9w5N/I6AExBzdvbQWVWGo3
rwtSLibQ7JcS/qHl24GLWrIUbgA9g6i6MkJLeQqrxsvXszNaMYKAPQpU4o+sStxexCzC2JX6Ywbw
RfSHTbh3mhEBT92X+y21v6AQBsbYKaJSGnfhbBJ8m3/7cudJcCYzCFtdOLsZSelzE+yG6q13cC5c
F380Wq8IT4HNCBm1dYB0AyS0MuBcZ2EX/W59EivAEpqk+K2IiQPIP4/zJj/TApI9H4kPQIX+NPOX
dgbUuMMO5DirtJ8tvOfhgnMSol06S0AAPW72diOrHG9eWs4ZfJZh5NCPlglOR7bzQPMtXXRSZbSO
W3FS0XORePzCa9ruyQ2Nl1SJTyDqpt5r7EtAAUBV1eEkR+zsAE6ZHD5y5LwY5d126uyIkYJl3BZE
RZ3XTvpIWP0mEf4O0zDFkNrz96UYKBumo7drAPWs3GtgyeFj/It2CW4MVBNxzvsJsdnoT4W8JTz+
/6SrISA7xzzUB1QHq076kXfFM8gbnY6FR4gTzCxY4Ljv19dOsogEH3qfZpUJG6h2CZALteXIWuo8
KAkLEyKbmx/SZGDeMOaXE2lrCqegkZAVZpshfWcdJKHCo+Z/TRH+y6Y/6QvFtX0yNNA5Vz+CkAn/
t1MpfZtHyYfR+hm15cJ9QS3e0mugimrjdy/yIBTqMNFUuPGjSmjaf+f/SrmnZjYsumsc6LFy4EEm
Y8AQSvZ4hBFsmS3FDry3wl3khkqAUq7CkUAkQUxLJFCuUvmLzIoCic8b1INrK5idXAiYlmU2uhY5
NVuH1Df4D63Ba7J/YvGDXNFrHCJYnULd9O9iyhZ59F4K2KLD+LErzH5YgHifEes0XGT4ubajA1gz
jzW9nqzIEuKL6bBUTos36HVmNcJKZE1nFDm0VPLGL3CmVn/t8p1u4VPjtNLYpYOLQfnXZLNJgfv5
kEiFZVzDewvWmjNJFwLqY9yH3E2TJsEQccUqnp0TPpu8L/0gNVQNoVYKymRfmRp0czr2BxIdv7qp
qXiZWRBXXUhfKbWjKIS1MNLoWI9+DpgmIrvq/ki5EwgWM+CBRsayAwsm7OhwzvwE8WjZsZNi/xvp
qoCXCpNiFrGBVmYvLsEgHAHxbJufhV3lEatJP0IWBmUqcN+HWsxK8xMLMOQwlTpRXqq5p9rkfdKk
5cIz90e7x3MTlHixdTnv/ErHmKRGeTXHekMFigsO9+Le7KCQeNP7mm0UyT5TwcmYvatFh7XjgcIr
db6OXpxPiqOUObHZrt77+NLpGcg0gCyaVJ0zJfRWQ8TSq4bWWtdr6VnepPo4X63Z0UzwyM9VTEu6
7Ei7rTb0qsw2wBGg+IZKXrYMnCTJNgDJk2Nw3rL1eQK3BRBB5rAysmv7Febk527x3za9ynRhg1sw
x3cpTbRHh919vcVKARdL44WvuI+UG5NkpxdvqRBTS5ew5kTNEL544KOjHV6CKrNPyiiH0XrAVa6U
k4MR/Fd0DMMWMeQ7SLLEfyeru1aQnp2baLDi5pOSGzmo5ueI7eKuf5uT9hyKRjNrirwrOx4FZsIe
Tc8dB70IpidhlkNYAS2LRhXeGt8khF27lG+YZyZVt/lZH1tzhzYvXQXbod0M8RboMbJMU3Z15MW0
uVINYpf5bPr/iJBEi6FtVRaSksKOnNljI6FdjStaRW9JqglNYQpGOaZuFXP8rJPUXJ3ad6VHupUx
KMsY/0Eat4UflXhFZ66V2A1dH4swyEzIDYfJTQx5jmqJZjS3SRNztSNNoHPQKzgxMCsRj5eI1H0H
tn1M8ClOcMPvzFGWCMSTW1e5/4RdzfxVG7EdT9JcvQy+1Ix8cRIf60AEy8aSEU1PGx48bx/1/IyT
LqwHVk/QaFH8uo8YBJBSuUO41CcvXO5xFFIq83P28/ztdzTHzWzJVO9VEIGZTTY4hHlFbnCzWmFv
oaJ61zEwaiBzqX1b7qgSXeof6Chcnr3o8O8gWJqGs5Dlo1ki6RDO5ND3gQ4f0j1XsrrFuYCXvu/S
KXtQEAEbw04JjWOvQyywRhSXBOe1HvYE3z6WwIXKAyF5yiYjiPdMclhBKVovH9t8nbrI50Z2ChV1
pYHIzh1pCuGwaEDUHI4haSJFy0g4hEHasbTLjb5870g4s9+kARRgN0EGk5sCrp0z3EfnxumWqDpO
KWECgBKeANKWcrLvwDZa066G7TuNwYyUosSf0Tud+xXmiMkh+5iAnZEWHuW1RDPqLGCrtaF+EwBe
SWj2MwCbTcjH4C9NzZql/cXywp1OYzoZcahfgkvOtHnYbyaN1/Zf+uefBSOYqTbbGbzcVRfJBeAk
0C8vdO26pPBEaWRruKIGgp21nbS0S2vZWd6WoiPrzPAPf3T/oaFwTKj5bggokdvZEnwuvreZwSGX
rHo9MFePH31GVsWgjCKgM+UATJgXTjyNaj9EKpksAxhIvyCEXfYs9XcRRUDiVFScPS3h17x4xmaf
AJbo09J7+bHyzihUQ9N8S7NdU6rBbsu+qeQfsFi2gbokHskxagY5C1zFunWiHs96YgrKQw5sG9oQ
WHhfuwpQoBuKttawI5T2FKM5aLHBF+CAUsd8jafqJByo86wASbrcPcgzRIGbZCak6S09B8ZHoBsL
A0ZLtZ23ivVUoOx623lDyxF0gCQAyF6KvjyavymtD2s7DE4c2bkAHPZvJhB1vf1Ztk3mKQcUqvNY
jUpAaIijTLTy0+3CvcoOfyDoVDZfYnvmp7unDy3vaaRrclCxLM/suppt31xO8Oiit8Q8GugN2m85
zazTN92Y0Nz3sd7DcsyACBEchu8rgBe6tzwRJjeko0hGyj2/S5J3yV37ILVdeasQ/OeUAtz3NvNs
l0O357nR76W+BFZlYej05HXvsPm4vd+bvzmziW2uPi0loqUOA06mzcWLprcfVczAqeSnt/raj55U
rjqgvf6BumMXtYinEYcH7EWExnoVqW2EaBmk5thpoaPW58XpiIYJ16Q1I6WQUnu8DCoF42XOHXX5
470z/q3pwjZ0IFxkd85eI0iboMB+andHGLpSDKrJFnNzPec0zMQtfidNwtqZR/UmDCGgunRoAqIN
QADGcW4WKTeSVDauVsEPzpC9XB49xbYGo0tQGg7dZqkLE4EpJhnppdK3AxxA3ORe4J8mzHhvJaLn
/EZyxPtLG2Knt7x9V4g+GeXGghCLBkXJmwse3Qw6eSXB55muVHYQc6Px9+d8HwFKEVKJFXdNbuEd
SkBPq7gVqWCa9WZ+g/1wUTuKLwBPlwX6hmCm8Opk5RZZOO+Y1iW7aZxqhPORvOFLw7Vzn8Vepka8
oN1ADFTcZEa7xdcZuZeWOGt+L8yLENeH0e9lhOmKXQEvGWKF5vKpKeF5JShm7P1x6tmCWh8Ss7YI
Oo7Mg/JgOS6n0bTLQbYxW/3mFd25057ERJ8GYsJTwjXZ+4VC868AtwqVMwBemeX5WLDhqrRfmrfs
lW32qG4AUuojKRk797LXNFMIriPKrygMjHVjsKXxAo8WKYyAysbFGGpEp6NpxpMomSH3qkftfdsR
Epp4gW/btfnZqu8HNgzBFs6UuqtxeCMSj7H1NuGOxF0iqVmpo3Sr3pbSCOVd41c99vDEo1GKZaLm
0YjDGqElkli6yP40b+RgY5dZrEzGs9y3zSSUIfJNuGGCORsQ6QEunmQeKSd03/TB8fGYSHmsNBjr
0eTqEH7SXMlA6kkTsehYIQfnn+qNm/AG+LnajHqSsn+qshN0HyUGFYCHlLsyem2oRZBQOPzZpU+7
+5mEUEGpFEk2BMhlYreAspSPkcXxwkuZDdaOra52GhvhY/GsTWyW+CsEC0mQaoDyQYl15xpgSZ8W
nXagTL1OOZNfj1QwG+iwl17m71JzO0nKp1MJ6jObJd3ZGEFSyBc+sGD1v7nVU/G5uUopc2rBpGyc
4Er3Fgctgn6BaceDvm6bWb526U4w6IqeAzOxOauH1E9efBV2yvTrXNwFZAkdQDeqerAhMUyUo1rI
NPOxboa/MlHoprL6I5xVb2R3ugOajeq5lrU6Je8xheHr3bUN4KAFITd+3p8BLS89FOkbCohmN9L1
R9mzRoNYGi5HaEKr6wrtdiwyXAtx8Ltik2W2EwXgcKARKW2cJlE2fF8XLhLWxVH9tBgZ0G8+MJ1K
uwO5gRVgv63tF7laBHmvYVovW6qqhgmeA+EPH0wnglpru2fvkYtqWbTe17m96FhlrDDp2bsrwNoQ
bmO/89YdP5tFANevtH0ox6mK3JxiRSbeiQcExuwXP3rKN4YD/dFV6/o/PS1TrHyHYA6V1jRlUl8m
l0VhMlm8fnEe87JvlghgWjFex7o3fmxMvuyi9xGnwS38ygqLHyxnF2Xc4UfaFU+H8ZzZsGbQsMvu
XB0GE/ibMyalo3ZwEOwGtf84HhUqwwj7sORfiT5jNFzCFN7vJ0FIEWyarNSHnMbJXLDyMjitCECI
3jTUtWISX+LUHoORcxwfYjCo9fmEwkTRxUNFqfhXeA6VOmINZPkzQqJXCTdbjH3AoXBQunL4FDSA
tlMoHoejPCRQwR0DE+q4Ruf/oTeOveVKed3EyGeorABkenpsBy6QYuc2w0BWm56+A6n6AnsIbv63
bGFQsr3SIhnNP/swa+SsELE0AyNsuhrAgmK59G6sdpI4WrzVk4aWG1pu0sz96GeoQJOidZjsCChx
EdztWGFS8b30LcBDIgk5xRBPsLsY4m7XWMg8fzH+JvaH5i3KnyIv1DnMLtBsKnzCVXzF2EfoMJD5
nhBFuXg6ca+IjHDfjvOkHD4eGCSVMhBMZkBLIYBiHvp/C4wMgltyWnbrGqjsXWpaBEcl33xNt/bT
zJgskvtL2YF5hTk85kdU0U7VgHuW2kaHEgGRsuWltIq22q6aE9F5J3t0Nnbss5SB3JIh89flz/NH
So8c+1wmbtwMu4Q6vyEijmkM1llIFcytuRc7ljj+7JHFBpjKsKBRK50vzmB/Fw/QWvNXthYBGYxy
XnCMnPgGwOhxmGWOiGlV1VQ67m0TVexn62buk68Ui2ntT6ieISVrdY7TQ7/rTy+/aVkRpvMfFpU+
oKoE6u17W7xuX+jDP8Jzwo7rKH9qE6b1Nf6Cgx6LNWIeZu3jOgOstXl/uXzkcU/2OSBJrtQkZAYU
Po1G8NfUrMtEteKfr7cWfpK6Mq77QaUP3p1cUJWx6GL1yUKP5ck0FpT8GXOZrMDkNOrp50GjQWHC
ub0qOGtXaM6LUziE4MKyPX9cgk2ny8+b4xqQ8OheWDPWBb4B1oze760YDu9nVCKy31/JJAwZ5Bgy
XxbVYVihA3ay43PsnL1CpiEWsP3FQf420nDskylMBmtPNE0kbAacnV2keq7Xn+oje8Pi4VxSB6Hf
iHSmOt2NRm3hxx2/nxsQFDYekfnHQSrpv7AijJ3O1HVc6SGPDA1VIbU2Ib1sJUmx3p8lwHBLEfWC
zVrTBrnQf/ActSYBYVsyH3nwnXSxdpiRnMepyDbkSeK2UHIUlbbfFMzYeBaMlTghiq7BDjQR7qAD
R5uckS1IVTiaOnoinv6AflIUDShZnLEllF2QfX7xKGJL0xya1FzAHTdUdB4yXvyJQswKWtn66FDJ
t/nDhOwkb9tNttOOtMd809hsruMl8uaEEa8nOOpzGCZYvKg3cxaZE8bfReFuq9udAAkdwW/ereoe
eZKERbWWy5ZxEl0dUQwEsFjU1SMs5cw1ZML4bT782MzukTQjEA1sn86DvN3pTWIE+U7nTPkOUt0G
YdEM0uFPyN2xgeiU8EM5yvQ+XsaQ1yKYUJk557AkJhW6+RWbbxfLpJ5i9doKdRWl41fKmouvRpSz
58XHACxfgtLS+KtuOM+9K3jlDbPV7yWkscGdxxBHaFNjrd+dr9Mw3aJmE69EOu+sJxwHlEH8n2Lw
ysuTARlol9qF8QEMgJpwJT49Z27Xjw2t9Ld03Ur4OsNtmWYtOmGOE2TP7R/ctnNI71d+Mt4Dt5Ai
lwFpawmZvBoDSvD2z++qRtUkPnReWGkJeQF0FoE52qxTB+Db9SOX7dZLU2ahXhu+nQGrFx6UVS4h
MbxElYZ5qWHFkf6P7nltPO0PYO4uUpdamRya0gshSBnT1FNVx1q+Tj6HfSCxEQ/7IZSQxFCrDBZ+
Auvio7zsqEcentaonItkn/eIk0lx/l1ZmYWySCN8vQIPuEYRlQCBY6D/IkeHsgtjo7SAAKkSdGyP
lxoiI/rbvCymF8S6OZEPhC6RZURi9xxj6hB95QKJDC0CdDiLNPRSHo8/b/2HRymj8R5bdXT94Njb
bBnhh8XlEOTDtlYN4vlig2FpKO/9mwApZ2e9rcLR1BUIpiC0JgRyAeF8sjSDtrMVZZycqNPlJKVm
0lMRrRYY38IT4kTPgn6MFdjHCD3un2DU4k51J0D/iknK4OPdW3JHZY5WEnaLRrZmRmREIYmHgm5g
6sVvd8R5847+5lNxRf5tUrdHeK3sBcoXlIQura62eY5FC5EoHhOv7uQ7W9UMAdeHPHITAtcInXrq
ulXnBCLFyXOi32wHeqjNR21TRj2QV9YHXuz/vpC1ggwEhDZsrel0Rlde1O9ZufiQycoLbeABpb78
kbDYZ3h43bAxEH4SUdqI/hDLsSvdhINt+3umo/w3A//swUY86VlK+pGZWv8D6F50IHP96yF2CmU1
zfKwO1oOMgri36hcyntPRQxv64zNNVvF/SDRuerBNP+VlyhOWdFsa+0wpoIqbcBfHH8s6cks5rVh
h5CNQ4zwhf+2aOHzVA/cqcLBNQJChyCxbOASNGWqn4qgiPOAJXTYManMm/pt82CruUiU71tC5mws
NCpcfVs8LSuijOlfZRgfsZPF4XuxprtcRvMdD6XYl05BA63mRnksjicz6TAX35LfilDfLACPoRdV
39ERghzbBm744h0rw+e/ovgVgrePtRnOCYWArY0+sX2o8Uva6l4hk5PfaZ+kiaFRoLlB3Xk9HbZG
dW/F7GkjUrkEFKPj6gJi3KmkZ/xbPpyhOWa913s3FJ1h9gZrr1ECdQ7w956oQcKz0G5MoM/EoiX1
QBPJ/Vilp9wgvvR6uMDjI0BVxJ7AGqa9XeBHpyXFqZ+O73rzd7cImG3F2OIVwzluNoJX4teywcqG
MWJ9Gs7+rsrX8M8HS/F7vt8rnBVY8ofbpu5Z2nJ68vObMUQrO2uV2dpJCWwq71kYcN4gNuWCKnto
1gnPV17W6eu/lvVVKD+j+Plosangb+rtFWbWbbuvpZ4RRS2QU2ZlX3L9v90RcIOSOYD9cyY3w9ST
+PNds56eB9FF3lzOyWu2h7gJqBjbcXiLQdLv1EOxICnmnw+YNt2765QB2aGDihgKsTYkx1bkDedd
iE/Su+unrjViFzGjtLlU3uJUoIEhiE26MA5DSN0ESxzWC3DPJxzi4WxWq1+HNnopuilztES65BkJ
ZzPz/F17tQGe7cYyWAELD6frX9GpoNxEyZuE446wqW/V5Afu0m+Teo2/pdzsMTER/4PL7ta/8kXQ
DieF6wKwz5wPZVyAbEp29CqcuMwEu5rPE8TFFMIoiUdpCgD0E6XnVDB56A1AenfWp8EM1n0Ic8AH
awOlVQV6OSvadwb9UGdXa22Vibf3kvp8fWcd0VWsIG50smxujPHF5lOLJVJW5vHoSpyWqdz5X8qr
wwdFJAD6jyKLgBDXQgCrtce/jnERgUD/GgFi1DbsJhNdBUrW0NdjVId5ErGEccWUe4aJ4oWHHZzU
FqoW/MXbaglQmD3XaWRBvb5jkvyPo50BxZE+ZXHqQdcj5r/GdAA5wnqbvTYSEG0zmih/R8ZKQRzP
gaALOfDgmqa+8bw98t6k83/ElAJ6XChr08e3Xg8TniW7xmNF8FO9i0NObhOvXHc411C4DDDBdP2M
URI/O3rL9I9vz4lgTNOAWWsYW+xetm/Vt4jcv41ypU5FC9yLvZTvazKREIZx1X0oNx3HGQfSx0v5
VhcZHwVgcXulMSVapbnkZcvyvX8tuV0mL/YVtZmR74hUFQeos8kuh5PD3ckCLMGyeyyGbcjvPeKZ
CHctyMzE796GJQIwnvFOcCw1JuqDpr1RcWfNm6Ju7tx0yQwtlBklbAe7jurt/Jsl5cFQX5h0dRju
rIwB0Rw/+OR7+VBx9R7YP8nnLe7csfuYMh0rmbDwpt0mwlYg/H++2A0iGKQZsYu6rVosAr1edghR
CdMI4XMlDo488ZSEc/lgOLFtl4OeSEeDo3xmIsitzkTIfsorYgku6iOKEyYTI2yHc3RtVfdmyVd8
WR5FH2KXKzutmcpJcxolOar0fRyH3yir8OlB6qqCIjIkRkr/eT7ihgKGuHFVbLN9F1Y6jGMRaV5b
ffz4wMpT0T5qkSTU0rD8lx9mb/KWOQdcaLDj1K9sJfHr7bfULBsBVSf7Ye4terqLG54P8wMkSj5F
lbkB9qP+xr9j1UEo+ztUWyWwAWXsarEAkXhjIiDBJB+VEllrcUHYfGluJ7nc1XnYRyhr5I9TLPVo
b1zCFnmuj66KKwBsDo1paRu6A+Qp/2EKB5grm+ScCm66wuM/mESqznbs/pwb+bfOFI1wwMaQYeMM
S/LwfZbGVS2aFQg0Wb01SL1L3OAKmGqjgqjsH0Lqhya5YeqycdBQj9lonMh2KpD0BjbnLcJ+V2f9
XYJGdakMZTi8x+0Z7e/x73O722iuo6tQ8JjltdpnwB2jNdz54onIPOjZxZTKNfHcsEH+IiMbhnGb
t3LE47bQ6v0iAJjwy6lWEMJGGL4CjdzNR7m1mzKry2z/yGFEUVNUDpNEG+N6OP2y2Bzfr+qz7LJF
m/jlcgp61Vj24aIk3TG6cg8ULMYVryTV9TqZwPqy64NuCyyxzi9xqkaiDcQKvLPklhQk9dz1oNpa
U9JUenNp+X81jGQq4K2K3+t1SUMX24So/pHXDSxXp+VITBBEmH0B7Hh6tG0scfFLSfyo14v+AqzT
o23Uz1V3o0ow0sXgfDHgm1WyWDO37oi2VkwN1v9DuWkmxPSSI7pdxHlViWHHupWEUxsHJx13zJjt
rgML9FGO69qsTgSRz5UwFucbNvYEJyNYBF3b9Mtc5+Jwkq3wFJ/mPN7eBNY3iLdMfoo+pnY+hi3v
CdQFw35s6Ko2CoK2UZhXVu8Hr4URDxGszhzUcRJoP/nrTd/tI+orBNmbRgrWIk6elnu582c5eh4U
oSrp3l+zlVndu61iKiyiB/u2+IoBOkVQHSHNHFJbIvxF55aYWaU2ReZwweE7kNb0Tm6jaMSme8R9
wRzARyuz02BSO4OP7b1NbOzmOoqqqXiudrMCOaefB5orNn8dn/Mdkr5lv3mr75V6RjLMmnU4m2y1
BUitWuuBS9slb7U2tDyeex3oKqcxR4Cuugk1ukmHhmpeiMgBnJZ6xe+JYIRlVWa7XZCFBNN5XpDM
szTy71pMyEiNPofMFFmH7KnZjcv8NejL2lLn5yIBrex1C6UiUDnk722CXuOH+BeQ3aTAlrKgB4FT
j3D37sOZmoX5njM4r0IZLQ2pWSfBBrHRB5ZBu4K1WjhLIY/gYO3nK2sJ8dPnNmwU+/AFLjeue/ZK
/3rehJInbGLwnZ61ScD/cB9TVJA4a/JeNASXUACtn7v84dYLYKu0G7fbL5JFuV+GeLlfwJY9NRrh
myA+3aLYABsY8TLk7L26DJ/q0Dwh9FZiXTGlB9cW4jx/qMunAFJZbUNloBLxKzJUHtyUvyR639tz
WsiD/nDba8i5f81mHolqp1G99HMTLRT/S6XuAUrlYvqOYjIpukpvuEImwcb/1RlO1E5+YWjChYKS
FJzWO5Cxw4rt9z5oRqUoBpbLDaIcwWQyhJF2z6HWIuWJkLeTmNx2NbS/5MuUIqQ+jEax1fxthgdX
z2hMlHeGqodBrLF9l3+/nG2M7m1nvZXSwoD4WI3PxZE6eL+v9kK2GLPWZaQAc9t3Ci3Ipn0x15UP
5VigLkESN76JQQUbVpY+iMW9z83bFK47EGZXakI+JUPsrYTzY18YH0rmr/1tlX5kf6+306+XTO8x
Om5nnXCqxebip5u1Hr4QNo52oEmwjCMQvHIcVV8Jrz5KZjk3V8BUejT/qfZZMbDyy53gW1GCq4la
yApE2zXgtZcN1D4EEEKmARDsph8rtpoc+49+ehuQOVHPuAXTZNNHLlLctUh3lWtaL6yIX6acoIAo
owtyHnxRvv0huM5mV44vobO5wkeEQcvUmtEvGWRY6ibMVoFq1adlZrypL6fgv0WsSmUO7k7r6nRZ
R2WyVD96D8XvDUeCZkL2zkm6s6U04Z2GjS6EGdwc9ULDgcuxM0kW0ITOxJYsg1lp0Bsb389VQoFK
zIgsZR4XdcBkucrPdiRze2l2bGhfj6CLy2Swb0A5e6McNhaweWzctUZ5Y3dyYScEij+FUKJlEoA5
3TU9IVSY/Ka7hlhaXHv2VlD5R/9G3WAphPGuMKmGeY7youCEMWmwwbChXMbdfXJg9Y4kZgsXJD9C
YbSK6mkf37QTUfHBUsJJyPqvatWSNPjz6RNV6OUHTohQS4cKd8dzfeoJwHpTm5s9iydxvkEEBnu/
mOTO7JvbbfDuBkaeebgdQU8zbDnqJKnE3FraZ4ATA1J2miLnkxSj8FP3FRmJJlcGnXAJHDAKOqmM
6YDVVg0FN0FD3Olhl2oE6o5bR3mZH412+CfUQaJlZX1WEGcoREL/2m0076IuY+p6ANT/zMLVpgJr
ndN5KbAQm5uH2IgQlUJ5HksD9BmlP1NHUUNT7wDXRKr/MY3kiMrCNFmpGm17GDnLgZp4UXIp112H
wSxnKj8mc18DsnFQuHkooyiazOkQcKuQbRNR2SD+kfi//4/IEoGmCYG7eXuCIOJTcZ1Pbm+3UT3p
EPlTr7F6W1DqAW/UwhsOZeSY1BV92iBkpx7C/Bg0uPol+/USBvfMmjwhg0Fj3/H5B8cGSBzN6gV2
R9fTWCPd8XNoOgRXeF93j9m4GhW91Gh2AdxrqzQq7ER2daINuwHZx2GNsZnzHou+YNl7XO+hOe4k
buYNju2YIC8SQhC2aP3jVkGF9oYI9ZScqMah7NGONueQOSGGfS8+RtvExqn3jKhSQ48maTEU0QA9
EjrzcSZrspmkju3hge6jgJ+yJjc53ZySUkrq9UBOSaRXb6W2P84b1KlfQ6g1vdpKuanjOlr5+HIo
PrC0ATzdjkTQ60A+WgLjSP+2DZKNROlmwF9nw4Ko955ZfjzEptczdgHrdgeec6dPR2s0PJ63jaVc
uMxeTTCKIKWqKiLBdwtI2NYPr5aVRjDML9nrzmgGFSEa21ScOTpxalLWMcPdA/WZF7TgOpXC2dSm
4WNK5HnS/Zv9AnGYXKd0xnMvbAnxUueW9z4VmtahQZog/7xmoHQrpcBc/5KGmZlnjDKspqLLdf5N
G2GW3TTm2TVsqvrnS3M7MzK6EjG1zSG8jEhO/5MsDmlX5sGpJTg8bkTmiTd2FVKAFpjE35dnytle
jri5+ODEwcPTsCtHjzTAb01GkqkZRPavBORwGfErrwabW1LBpv7gd/BHtWFy0si1bjoISmLyQp3R
JXVxR6f8aRDXudAS/znHaWk50ISZVAtVJE6vJacEovJNNHYcS5+s+q0phNg2cbo9Z3lWYjrta6jH
xyxc72grkgFeDg0/nPhKvyxSezhsDRUIhTqkAPeWPnrS69dcXotXFAmaW105hmewtcXt5my32SJl
xL39fAiS7Wee0Wzq2sJSHs98S/81CktQJBJsl7tQog1cGwo8s7+NKdIGMyl41Dyyywp+VdUFZS6r
tTVznxz7jos6mTBhSvt2kLxOF3bJEFTxrO+Sdv9BLvAY0VCymLky0+kqvuhUC+lh2U5x55XiOSG9
goNbzTVG3Fpr0+4vmkYxDassXTPTFKQRch4I+8P7Nk8q3OjJWdZQY2fpwAWoOXosPTZ9bT6Y0tjJ
oTpFa3f/7W1RaNozSO30/RhPYHcPf+5IpxGGfquMaWBhuM/ShwFx7E85pAvmUoIjVDefSZ1WvuIH
R3h9TOwZD6TDWqyBHo6xrvsK2TLj5afOrxXpuJgZPQkQXqmxMNKTeRn1bp/s4Ba3XBCPSFtHEmnZ
lWn/sZEzNskGSJ2lh9bivo5jKmxsIypaQr4AbvU3+2gQH+t32hEFB6LP1Pv9Z+ixAT8yA2FU4RmN
Jir7JAxsGcJwbFg+b5dQXjoaQ/eiIN8d9bFlenpFjBckyt4UH06KK1kf7Agm/rVvBmhhmwv46BL/
l50awkXFIJHw6a9zgfRKowoqCEZ9eh/2K03QQZnNauX/wXAAuUltB5K88DUE/dXwVDze1tNSom6A
ZN3BEzWNXupdh7kbkD0Q3Kk9+Tmdw3pHZHrZKFx5NkM4sLFxuKyjyhffO1gRKCKPbO9B83L+Aq+9
T2eZWSldqdi704TXlb+MoOeJ8lHWsKP7yZ8NMT5Klyq6iKL15Ry5k45OMNWv/WOilJt2DbT2gePo
fVVVEeyWakiwM4Y3qDAuDz0V1FIlOdDLZi8xApWejpllw+EgyHAKIeRE4F4YfqeWXHrTOOH+prAF
mbZcWe+sZ4jt4MpnI2A5W2iS4QkimgBA/5MBbxEOdQlaEwrbGsV1H37dan71Ur1l3ZrO93/EEYD1
7RDCHhsP1ccVzUhor120aEAwXWQcsLwFEg0oB3VTAnjUjiDOh8zBUJc6nFCuiaZjqmqwEe7+Dsoq
YKpGPeHt7QIKibQUoydyBQhBch0+HIz4Y5Ve4UtLtKSF98wTe5FlUrqx+cIOPcz1Gew8mqOoKhby
7QlNTdJ2JhJjo/CQ46TVuCihdXooZVqFyzc63e82gkRmzBAFOTjVxYkXs2fKuamrFdz+0NcldOsH
SeI5LdPmEqIEkmWuHWTGOxCVG/Swg/ax7+Pc5D0jPzBDOECobd6Eum0l6LFwSuzG+sES0fV4wSQt
Uz9j/QA67VQf005DiKrqOe2cQgSRPbuFs9QlEKxD3vmQzNT1oCwPHZ14i73a0H8X6yZtbHwnQmNS
fLQyeO+ERpU+H5pp6o8MpaDK/tuhUyCTQj10GaiJlCPpc+AHcL50Mss4Izu2mrg3D9vlEk7PvYrg
wJnKOO9SZchUrN0QoWu/GQaSF6pn1hVlXOjYvRa42x/0GrCWmpg1lx4GODlYO8JK/EbtPUuSYtCR
gLrnoDSTs2zx1hy4K4eiB+EvWPBKoVqcBxLuO2cm+uZpnFCR2UJngQo9zPP0pEQUwfA0jVGTrS6W
9cDEfGIWsR3gmWiieH6XhC60NIKSGpVjCZ5OiPIRQ+J83Kp00j0JvmB88CR8lKZo3dACt1t0X+5N
03auPs+MWJy/qNBKR6E9150qDWoVoKGTqvro1dZ5DqJQfF77oQKxunJRqsU9wzycQdmlJjTE9Mhk
F71Bcq3AHXTQwZERLOUgZMg5gbRmz6jTl/nxJ4kVtrP5JS7v0jESbMUVtqnzXULk2bANu4EPQV3A
Emn7hiwoV55+OrTbCUd7VNsIPB2JvJcIHHWN4OWuuvBoWaTqZLgF1M89bFIsj5oi6TXTrTVcg0d+
2mDQ6Tc6rWOiuMoGL+9xMQ6d6TihtJZWKvyWQXe0NAQF+cc7RpD15Kvxu9HGBBSfkJTqzwK7K/2c
8Yr7um6kEkA67wvbvNiUpm9O/e/i1guhjJV6KyrhPGYb3dM8do1WcN1nvFLHA5NYH9D+0ZEnBo5k
8/LZGw+T8q9peTITeUv6YPepcmLyqid5a98YEPBQxI9aYTwO41iG1OTXWlXlZ9nAYuJ3nh+vr62n
1rrw4RTlHmslS4F0ZsDm2zyPV4IXJyTfB8Aoj8QXFZ2Gv843NHKw7x4TPr3rvBnUx8g8oBQ6FSEA
q0LrcfVgTIH6amNNVsUOof86IRHdimmrzlmomccFJMZk4uDODY3q+bfrJuwLLJVxQCcKhObI50wy
4cHtAXoA2pTcSuweH63yJM4GTGMtYMLZ7CKY+MsRwWt21ImvpOkdwKyCyxCGGnEAxiw5RODyOtlT
7q7pO/FI85K9ZqgWQLOGUp4tRMaET5l998P+mT0i2FS/RNthYQvwIhnNX+8VW4BoqL2UPlZzbnUS
VynHWNz+pOapaI8If7FoSq5gMoyx6I7QF+xdj5pm8jo4h8G1Za2JAA0iR2fx2ZmS7oc/D7+CwlfH
2P4KYxlfmlMpc/Hjecb7DAJXc6QcFREfFuIGYbn6U4VguD6SHPntRBDI8liBSNAj06VsaUEKAJLO
OeM1qSjw/X1mEz1K/L/T4dxm1cUa6zqJ3480LfcG6uLU4shGIEBMNR5Vrdn15Z47OemVOXTS3/w5
DHj1BIEFjZh1EDV+vV/zzqHY2VwQD87fE+k32rXOzYJiSG4uEPF8+HtckjyohwoRF2PyiqnnWsgg
qFYliA5XDXjiljAZs+BW7eGFYq2dg2h2CwTOY23Q9oKiujR/JsQwyPn1PH6x6i8uVEcCXSllOx/j
/suYa88D8ugeINLEAp4cqh2hrRB2HinZ5xhBy567lCy2GKQtrMEhQIcjLL+RP06r56cXoCju6b0E
XtBf4fCS1z9uJtooZ68uqsrwxDd1ZSqHX/fLdA7RPQ2VctSQHi+Q/nzv7pGVZm61gb/c++kLp/Cr
zuG7E2wtFY6Vt2zZYNzxsh5QKdwnlFAn5mvtiK24FrtxRK9/gn7WjN2YwjjPGXjuUJ7IfDPcQvOE
DWYtFM0UY4H5U/iaza6/lCBcsMs9LZRsvCzsBHMmSzVWKRKptTR0PgsBAk0YGVYHrC6X7vrn9RTJ
g98kakmINh9OD1MiyIi9XajgqrUCyT0IxtU5MQmgdGG+POKvm1pDsGhN74g1jzzk2K+iOJ56EtXw
FPcUNSeZTyWVN/+2BWHYg43SCkCSW+oLkcLyFQL6s4yDHv4ibGYh2AIZlcZtjch5D4QGUIm4tD+X
Eocui4Xsfg+I1KwiXKfqRdftCnEHfNukoRQjju0+i67RE53/1ZEWKHxitcHMFXQgkoEBPnOrNA7o
XGi8qQn8sfWtDe1mYhMVSxfjIDRanX/hgy0bA3SYkBFlmsD54rEzPJ7IqWZKE3UhnucXB3dLOQvv
hwn2YoPKKA6bLIqFZopZGlcYAnJZSMI9cEwnKpIuK6M0GTSy7iSSV02I1IJ+q7k0Fabry/5s1zRg
Q31zGsr4WHAGVSRwsZsvDY8DNKUHhg9CgqelpNT5HDNimKFaXXC+YjNZ1LZXyIEKiZNp8bd9WlIS
P1P4kBjbZnewK1TRLRWhRsCqTsMd2iYybyQ6WwqzpnSEKsy+7LM0zj6t/qk+iuzv9vasXtnwPrsg
yEhSull8XaFzYz70V51mxWiARiqFPGExpn/hEwph+Zow5VG1YJhAeIYWZTSLejTsxLJ5av8XkETi
42+tBkJ+QlDLS13iv1fd1E8kA7dBTf1GNv5EWokQxCGEyshC0D8Ul7ztEYo903KfWR9CNcC8X/qv
23IjYNnase2T7C7gXxz4Tqz3Hlxsbju/rJu9nSDJ3IB56JaFbCWKdWd9o9oDB0ehmrYGmQna8PTy
7QKxHubxakjTdW+CdNIuBmXHGHy4w8DOzYZlAKAY/MN+yilYqe3Gq3LmEeT4/iE+01AQp9qLYMol
tRP/P/bVk4O7VEczOFmeXxTOeSnEEtNSf/vN7nrDjL04KF3Ybc9W1gf905qdZSSRfdubxIgIkHMr
iC58x9XT2gU8dA8DdurTIXVs5kpQEZFrUKzB+JKqb7/WdPdX+rozr81Fi4z/qSIDS4ru/+z9Oiwr
1wNmQflgChwd+W7LF4rZQgeGKIoxI87oSU4duMuajgIxLDQVffiaCPTDXPBSwyll+bQ3BCDDucbM
99qs4AChKs4f2ljETYvhwSLSkfnToPfhPhI2ozICzebsatmQBjpBGsVwW1RWp1oxf7oBfWx139XP
7xsoY2U7XNWxAmxefxXD3ftEKoMR7qD8VhfyrfiIfKIjWE8h6gizGKgnzg/irpTa1XnHFAfXZGHZ
Rqr4e5v7+A18JQwQeT/lttaQ4aJKAYuhkp9DJbaez2UoGeeqtCXmvJpfLm8UXH67gXbtyZbIaxUU
K8ECu49pvt0er04R9Tc6oCCzXlfEPBuQfkWkRzetpzMtkn6XBLkqQIbFcURsO1BkdhP9OTc4oN1v
kJ5qDM1ik8zwkbvKd0NB0VQNVV0vPb8wVhw6K79X/P6Q5sAnO6h5e8ql4qWL3N46kiwBsdsoPk4s
/cSSuQRXSfEcxMxfqmL4LtuWjLYK7LsxXUOtLJYeMeCvvIuM1BtgWnpqwc/e9Ym3SiWFy80Q8Fes
E4FwVClKMckLgLyWPRPjT8dHnFVlBf3+jzgKQeCkgmWDpvW5AepYD9a2VJjJsNi2hnrQv8yl+Uec
9rUtpzPyXPlWC9B+1X6yWJ4T6TvNqE5KUPc6JX+EgXhm4di9XD9XD3Lg+Kg5ZrONYcTYYtlzgrc2
NvGIhj1F1hpgMmjI0ydpnYz7af9jOQe58+ADrVACqLNemDs4sOptAF2RtL928fTRTlaIeQ9GYA7T
kBDTa01kO7c5CbOraBjM+LGGN0lGGfdk/MrezfVW4CPrlPxsmo81dkbBncCt+DZCqrRYNypvQ1D8
5nhp1mrL6mB1QuFaxabSI347SCR7daUwCXWqetcJQ1j+TCa4ct8HI2wIi9e7IjL2h36zDeCVyU84
QQlduSRL9FUGlWYoDxSJlxz9BL7uKG01Ecs5i8F80h2hJ+ZGqAzEGntC6MkS77WdJsC1A2HHcE+s
PncoMH59XdEcJxe1gZ4bY11O58n+l/gj78Cw9xN1YydM88472XpvdwwCLKlFJ4ST+L1jPwStW4h5
sQbFUiQ3cZcxpcXifQtwW4cDgr8wob9YpTJZGOmiH7X5ZjgEECE1K7Of2u1JGlpgRcaEslUjAbPt
fl2SYYrAXlTtvKUn+1FyMzY7PhqjKx1hgW9+AiyUrJJcJsQp6FSKDS+iIC+cYSPn8pIRTYyc3lyw
KqGrGSsBWKiujdF+fDFtqsFKQz73M7nOrmS7XXlADNRW5XlsFUO/koje7f/yQhPdJ63xKVRIZwLd
spktr+3n/aP85EZ3lyEsprR9TT/CESqcHmxoN+mfpu6+grOe6edu/StMSZocTFjvO9t21m8JBfKd
mUMNfJ5UXYnrUb9GafzaYhgG1aMjoliRVhKuqlF8GVMrBWpp34j0RqapWn9dyg8+6EsFqSUuTKL8
1FVBnRR44CddeE2Zzg9Fuhp64W0nMToEl9mvW4MWdfpr6lIGBOwBplx4o3dQoZPLxtQjlmfygnQA
6X7HQfJsDUONSn2zbxBpulpRyxTAMFGFAQHMtp+MpVOBGIyVGsXJHgW7tq9UBMEklXyyB112YpJk
dU21PBITO0udzoK3FFEQ9ROqo0uBDvDfmSQCJLmSkkP/SYvJJQQsDdwRmz9LjWXHeXVwcpc5Vwx6
uTuK49qqnJ+YCnHHlVJDfgVFb8CF/tzdjVO5ULzTI7/3aW16US/RYGTPBN08vUprYYCV6NT0Rft3
j/n6Q8NTIqc40LtG3/67YQY1pzaQZbG570xTzOSfzweXgF2rciLW5AgLINzPIPRMPWbeMQJZYbV9
W2ph4gCvo6+XR+OhOKgALXrt8VIqv9+dAvX5RSfSKmMx7WK3nW5m9jVLxFh667/y/SGmuCDkTig0
LgxV7gWCkw3Z6f4CGUEB4UK7HyJlxBb8p7RC2yIqTnORDyfasggcwosRU6dRQYClLqcUqJxQsMfY
3hDRq8vrXHSfar36+KopHOJUFWyi19pKCLijXJPyj4kYv9qZBspw1kHduGE8YBvsq98se7udpeH0
AwbRSSexDTv/aPAhhOt8sq2rIXEFbqJe/ZOkg4uqQOBbiBMWypCb0lIu2jGvoTn5MmYi/b71Ozmi
dH3qrQr64zJvbGG0mr5MsLTESoqnX1hVaegPSHM24J4Fypr3PbOaHfpWMdX/c1V/fS0jes7MyZey
zdIUHXZVgDVbM1Qt+nHkg+p/8MOadxlb5lNro5AKEWOJMuYuxhxQz772+alyi5eAE4iMG9U/Oa+u
L9l3/qF5PiKBWBlPkh+AJKpnYZjJW/VWpvosxFjRsFa1x+OdEdpBd273KQw4tUqi6f8s6MV1hhbb
Va55HQbi5w5E9NlTB9jPUpkERSW2PueNwpffifRDBs3vQ+C+uxECP/S5CpikOFXDdFJUnMIwORlP
NGSZrRAu5Kp1jRGL0wd+pV0cH+RHIaIvnyTBV8wNCByjHsoO37QVW9hB/P++VOxO4FRIMr0yqkQb
rQjsJGcAKOeFmKoy4AszGNdfB/mWQbNrv1X/ajcH+9OpL1AIqf//2VlLfakvBDjXHUS5Ty4L90Zy
BEeMKamxq7Db497KpSC92Q89/MBEeUrf0IbvM/U+K+BFaQXCU1VZqjIWz+GIkqOdgamC3K7N58D6
WgOcLVcvZA81YP9ypelbNY/1eekVtKaQyvpOjva63j88YaOcUT27XClkJREtf5twvA/rXoZXOhqY
XD0bvzh+K7hyL0l8lPR+qcG55XiWOd7YtWhSshNJVZT4KA4MbIXFTf5HMadi/4AW9CoMSsiHh2eC
fusGfdbT/YxyDI5ah0ahH1W8tpyonWDwmhkHaGHmRodw+gehcOyhE66Sa8wqiADsflPctDqx7BrF
+P/x5ihAWM8i/Wkbf9SYBnoGbhNAscNWLsAh2XFgDm3i77xCp4upJCrCbvf7uPu2/M5TraUJOWfX
AvfNGd6MCHOY6IOl2iwjdgG/JJ46FYGoAOJY7QHZZouGn1tjz3uspaEoawcWtA8lmjeIF7197E+y
6y0PU4RpqHg4lOeyq9ulWAS6xf9Fgz+VBi5EyXv+F3TaAjZ16xNnkPrReQSTVc2AFg7zs2Ta+WyI
ZFAZb+XRG0xJ4yUSjorlN5BhEGQzoY3riH/eXqwzwz15+m/YQIdxRM0JkLLJr8qUdrp/vvYU5+Gr
T+pR9G4CNVCb3RpU5a3Zl6X/lREL2/PLu8M6kgQ6kk/tqBWgcSdsBqz5fwG7NbgxVaY+4qUyLjnx
jcKiON2sAENYwJQl3vx9cNc9SkATk9JdgRXK4n2CRvfdpcCt4WgHAwaDTrHbAOmryc1Hl4gVfCO1
5mkqil4aBg5rWJ0ny7vSSvHdvGWFBAYTCtxWOWXJNd2E32WAXyC8TEjSp32rPgjXYmu/STd9X6Rl
BIST0Fs7xxW5WNPdT8Lkhq20u2jH0UegOBirY+AKVJZGli7QGYRHa/BoTEJImIR9EPl17gAXXHfm
ARH9SbUMbYe3stbKGtqM7kbKfghR2eFehADQsHqzkA67Pt+/BYXeM7X0vLIdINbYZTzq0Nv6crwV
mptoUC7iqr0MpkHA/QQGqvObuS76EAII1OLYUyH9Eyq/netEJJiPYqRh0nCfUbS0NG9QUhv0qAre
wT/toqEREz+Bugat6zLWPWIo+i+AXdhRVz6v4lbM8xfIN7FOqbZ4stATtbKGOGcqswKAb8uU9sRQ
dyyPWXI7DFztp0Rz3WeAtk6sG5a9e0z0aTg36lKsgjhB5ZIVZboiX3gNc2oPFIh/tF/O/yAaYoqf
dpR+J59XWnAF3gD10/SfHtw2X5Y2R6lP7ASssYj5jOEuIzXpEdPnehWcRdjyee07wXf2HFcAjSNt
MqdrPyX7gp6fszCwgmhfuWzdV8vcAty0YB8FbMt5/lZJWUIaW1KA/NwQ/vPAqU1fB0HrOqg5Y+hc
9Omt3EYDjK46KiBbgIDU9AEwRzTZmj/7qHd7THZ/culJhGg+OMtVocHPPkhKfk07fF2zt4cGucFM
DWEIrvpCY+OiUSx1XCNx6IhEH39P2VwK0E83sO3unDVyRbVOu/jyvTSOd3Z4E1q1eKZSP4bj+vJL
QDYFqbcCwOTs84xYQLxN/IdeRQVqUFybX3ngDUS4oHZOHIJUWU7MeU5dcT7wmrPkCxX7KLkP7jgp
ZAuKl9zdP+Az8CkW8uGf+M7WWrUcbyD9NbEqAAdcUR4O7IS/OLm5NAcdJvmHiengAoF+XdfcAhuT
gHy/wPZNGCFp4aBc045XbWlFE+zh5CQgCKrTbn6hmu257xcckdXCEIQUpWYA1+Pt0xdiOQyVyPsw
LUMA05V3jDspr6ZToFYFEhaD0JQVitj13lGZqLM4yXsEPLLwDDUGfviqmODjA+jFS7f+tRT3k1lA
txXE6sMKB2mU6jlWHM1uie3CeJZJtwbR/rjQDF1zT/ARDyMRQ1yH2Z9VQ3RJrBz6qqy17THG7WYT
BZKVo2ezmWu7rRXTAv2Oht5xxPKNYfRlOZlIg4jtWUscVfuNla7EroUOQhhrxvUKqRw0qfGqq2lz
NsWSTOqFa4F2u0QRhhc+haSC10A4a4kSz+RMrm3lZcXyWg5siSIZ3q3TSYMKoXgXLgsOYHesvCtw
3+7xiK6MkvjHoSw9sWXysY3T8dm+DfcN0j0Y1LVrLKLssVKgh0Ph5MC31AIovBJmcdTm6vkssC3w
GGFtOcyQ1zwPeJIGXd8eKagl61nJJXPZR8eslvid9jnavQa6L8Z5Zr3KYe1rj9FqsEhbeM7pOzOA
LrKZAgZqqEndXaYdbC2N6wd9U3a9Z1pN7CBBlQm9NIhoPU72YkaZ+0ihWjLBqByaiOG9zbtx2m6j
cSnIiJbdq/mSGnp5i0+H6XiBQatCnYd5BwnF6ypySgPgEqpI1Ch+eO11zQ+l24nibrxD2JNN/Za4
O19UNuL9te8pZ2KX0OR2yWT/9vYxDAShdDc8Q4VC1WhXaHPb/6+fy3vQA/n9rwh/VEWaen9M2o4z
SlzDLaDqQV1reDqie/flYgj7YR432ls9gP+niNrvXw0a11TMUmDsPmtyHl5gXOlO92j7RTbOWiLw
qs6bR+z+J1Booj8QAZ0UmvUHMpHh3UfTty/OlHgoQIirwTHTzFt/7VhH6AR8f9GKdrQAq1AmgFQ3
pmnNSsWJIXlQ8Y3co9hEpLpB0GpX7qXOnwJaSui4CUSmJlIQeXUPJ9xlUpg1L/7HmpyrjkbnexnX
D5Ln8BnjzhusuiYPrrMAVfI2nLZfpiJ1jN6yKbVcX5iEFla8eM5erK7JTi3qiV8EZoipAZarrulc
MyOSZ8EPeB6pDd3iEhEA0YAvb1QcIcRIQOo4TFqRBo6SVEkYd/XKjJ0LpI5XoX82vzGw189eM3GL
bXJ9Qo0YU5jIl/kmo3jGOeK7u2E3KpQcr9YzZ54FX6A2aOhgn+CxMAZqvNujQLfMy+SwEfOIuhXu
Cv3BraROsenER24eMcwb4jAbKiclNkiW8Gm7qSwAcV85LCDL+7e0PdxcSrgZEnlHjNLqnvtFJOYo
9TW5y93Y8Kpvf/AX8uPOn744zJNxK9ft+D7Ip4F58/pzZjEOUWzraDwqHSlsMDH7zktEs2go14Dg
W369iCe762upsAgQnssJHBoUlJViFR9jE65CEir+0DUCcD0Zrk/9SMDIOJhVNe584JTYzjNlr8RH
KkdtFOjewJ/IVI5KjSY4lDMaauW9T53uiZeRcjmp9TwGYOOigvoQVe4NIO+J2iemwQtmnxL8LbbM
BS3JuAgm1aY2QQ/haXTARRdwZBpddnPlXF/K8tcRXY+BmkzIpklF1oau3ow7P0AE5WM68vYzsJom
t4kjmReBFL0x3Qs1tZgv31VMEGEVeM5zu556UhTiseYU6sVbCKV4FX0Zgo9WsDH1+sxyuMByk69Y
fzLsRiVcTUKUIbZFKt3bHK+2JoyDSZYc21JXjeJLjUR6DjcLb5Jh2MHtysKiWmZtJqu9R36nQ7Cf
ZeTBSHgSxFw/3DCY8y/72ggQqv1aKJUz2/w+hdpFcOtnjXeHWj2jayJ/HoCkeB7hvtcovJ4Qi+4U
5EO7GIfuZJX2bSBax7AOxKVHjUThPMj2Y1jgai/etGaUbAKmtk7EIvIZOdaxiot7PWWgSBxgOtes
Y40n01FOOK9SU15S//T09kSAr1mTQjBPsxXRgnjO0FG1su4d2n1YHPBQg2INeQrxu+LD6ktfHsr2
Cc0PswRbv/qQTSrq2dmWpG4AfMj4C6DQNU08Q07+0+Q4p3WkdL3XlTcb8aVnn1Dc/91QlO0/7fT+
i3WmdYx5cuDb63t0sZsT0a4NcSaycB8baJ9SMKwL/sar48WdOylREhcnHRrKoZn9Ys/DhSzl4078
rT3HtzfulxJzXFQMRwSh+wn8VXPfkO9XRBA6quKWZ/pwkVsHvudOBSx/5yHPhIr3H4G7/hUdjVO6
aph1j/5dHOZWQzO7S0YhcJcbA01Cemscn5G+7RycxOy623dtZesYfMZ1rWWiwrIFQgFpTz+ga3LM
Q9te7AZUQvuUgM77kvgMbj1pK79XnKFDyh9GGf0/FMeVTbmycBXq66LoVqwfMiQUmdANVvimj2zt
H2tKTN5FfHrPhfTV6RW7paM+m8/vgC9ik9rk+QPeKYwqYlnPDPcuhY/oTizmcY3mXyHRQJGyLSvw
UPmxmQhD2BX92qA9+39nKs2P3DVWnKh8EmKp4ZO0QmRn+FnhDAYYOrDSOgHLdcQmAruUJVY7pP0A
02FGhUbW52tnmE1vdrUXaXwM8XAlz3fYE7jRn+zAZHVvaCtFKvw8dGGtAlkYYl6t8d60j3Khhexq
EVdhaGeDHKWQEBzVkXseISdLgZYkLTqgsSKQ1Q6XKec0hR9yJc+xzgIFDzBOnGmZsPbJJvjWU4vI
cKNUJ6klEDxR+O4n+FMcOW05lKnPYHJcfK6bnZQPq4vlq+im2UQ1jrl2e6DKvL+LVG4uWTu2Ld0K
qnyhH2jEpwn84NIzWW+sUnkrO1hXCBxU+DtreG6iOr0N0TiUnHNhho5kRTxoGOV0e97RdfLYwj+k
NAZBSxAgGUR+b/c9zjwLdYpk1oUd0xWnXJOV1e2osIAN8aYubDtgBQZsOnqgNX37v2fnwUWbe9Sy
br2I8SHnOdW3ye9fVVb+rUdOV+GMRQwRy9wYwojjw9YpxspVwsfKOb8y1zrpfrCKu4U16BFd/wpD
qEo6mMkBrb+psp6WjZjtDscccRdGEYGaDKRjl68vcwADbZrZc87ZJOCzajeiGfSXPOqhkzZAmlwK
n8J/t03vF20LW0u83h6jZY6EoW3UtmfVfAnkle//YENo8cbnblRI3omylISeHOCRn+kLj7mbuKjj
tZgc0+Z54Ees7r5xXte4sqnyunQ3lBNY/Y9MsIxpp1Jwc7X1DYKrI7XnY/ruqFKtRghPtzjPdx5t
RkEHor/64e8fW/N+e80Vemxvd3N3zLzOYZPtK5xuWwlVIB8dOIFE+oWe7Qrt0AfSHBDtdYVjqhNQ
mrFoU6eHx7ptSDEIaIX5vd3LcNJsx+mwxK5PGz7gaEuMOpkarzQyjHxxqRG0eo7Vh0lrCbKjjy5j
0K+1H5Xgv2NfHo7T0Y1NcYpXu7J3oX6iqxA3eClQWlQEm6/tKbEW1M5S8eNuBmV4glRrRx3nyLNa
rtxuMTY+G7j3Y7S55pKgM8HedH3YwXuuhEo/3opK0pDj+QY9YeiqXgpRnA48dCVsx2us4YkfLr1R
48JL6hMhR9xCFQbDUZX/Ly6cSGxeKRGmkvy7opqtWi3WkbfHnVEZ/rbt973SrMgJy4bxtRKscoBQ
aBIsCCG/wTGeukR3Dk3lJnvSHmlpbUnKiBAZhDET9OitKUnJMHJmeIYUmTjZ5cmMCPc70W2br0JC
FnbToj2hGkvUFcKGza91iAx+hb0/+4Lu3O6Q/LlQiM8If9dJoP1M+1ibaJt/MZx5b97zwlTxcdLR
a6s0FDZC8/RUsjdzntryoUrf4BZKKxKedSh9PGPKiQJnos0Z/4db4xvAaKCVvdgkVacpeZOBxnOy
sINWua21/Do5QVvHGFTB0BgmDx476cxCSghH8+lLYBnmrfypXSxkwvnuFItXPPy831LlgvHK/c+3
/niWEgTf+jzLmkGqo3VLHLbVjtRH2cLFRFOta+/tjh3/gvwdtt7q0Oy+jalqVpVuY2XfxRUyg75R
pdwINy+Hue9SvX/XZBzGpf+eU26FOITSxNo0tyWDvFIVvnP8TF8RPstai8uxczU6+fUFkJj2I2qz
vYp9iXJA5kqdPg6DE7YlmBc4afFh1gyONrxUs0FCXYXlynjnCASVK/vXZ8RYJP6C4qyCUGWoGMzS
LZXMqrVcy4rvP/zmrocIEpJOR+WmRrg6tS1AF6SvCDmRrImrZwA/sbLB1o5paaQJh3aAzq2CV/uZ
+dHW/K/6fSNwRV05rtKq/q/1HKkTGEQcuQTe4NaFBVWGknUtjxKBn7iuRMoSUA87rv3xwa0bPcoG
5W3L4mKFlEYFH+sylwgesCr0QI1Jn9qo6R9BdG+Eyir+AtAJbbiM+IhLiQ3ROcXxTm57lZqjLB1U
uavzdDuMgvKGdQam+Pn0J773gs3cdRZR0zgM74OIhEoI3jsgBFFUJNe/B1208fBi37v+VstwrzrD
AW1KNPZ3jNxxVOu7smDWY+uQvIZ+QChgYnhU+cd867yHeNzjkAwyN4KTipb1CKgjdQUCjCP+f87V
1TfEqfhI34MrwGcVn4auhhT5eaT+e8qNR54GYzchHxc3efGYH/EewKQeyqw8ndEL8NFp40Us84tq
SUkt7Hz60T8xH5eiKhiq3TRF8LGsj/MRu4m3ps1Ui4FKdhCmENf+AAhnJaOCGWh81lFAYJ18HdGy
45fcm872xSHngk38mf/Taph+oMoIvq8WvJa/YMIzSGFuclQrWTknScoGi3UdKi95Epp8rX/JgMn1
wRYtnjJoL6f73sDlNRp9G5/zDME/RGOQsAds8bGzUwFZDC1GbFR3dpU2eXGcJUg0G3dGJnNbHo0n
K/l/Ov08hhrJUhsSyv9ILkSUM2aeZxcg95P0rU/P7sYIZmf4f2Yd9hSBUdvkQeR+bdpc8PsIg4GM
K8A28GeS4ZOxWB51lKzPvLuaQ53eO5mrOAxcN+LtGM8SSopUioirNdgDuB/3r/ctsfjNqSdH5H3b
NUAaKRR15qkQiJwt6ijmZiqPRRCMFiI5TDlIxSzlHoscn1TQz+9+4SuhAVS6AV+N06mS7KCPPjGO
ne51tt7CUhkwYMwCNxr0iYCXh/YXegjPEhD+x0MXNBBTQImZ8zHeCdcIwyx9vPmC3a+Q9bvI+QXi
/A+urcAUMo5DnZOEBtV7H3SWYJMVksn739197lazDyo7MH/hp3qVA4qoktcX5axykXHeP8VHoK29
1IfhmrhrzO45n9iINoj12h/eQ1OVEdZ3eEFJy3+hVRmsBxkw4oChftj2YJ/IdWiHArx27sjecSaW
un8VO/mRXuz6r321Pst586p5NIBgABPn+25SpCxDhLVOAdJ3MKp5fb3g67vs7OHdau4irMaqcWPD
HgV7cHVd3Eb9DalaNnhnct+Q/ZiX/7VEzezXK68ErDuzU5pDmKJKF29d58S4gVVi1XoB55s/eSEf
t9UcXmWjj2TuSLZJSgoQ6e+7gqy6sc1dIdJXw/7SC0x5ChfhCuxKPqNmZR+Mb3sIHDr6ls5FKF9q
2oy9pI9nUNahBVF2S9385msHlfrZcrv4qAZ+DFDzZpIsPH6zJIADNF1whpzc3XmvukkioLWk81Vt
LVsHESZ2TGwyTPRHsxrnXlKoBIVNffQ+IXQcbsUmr3Mz7LANWtMi66rKvyhcCHVh6JVMfvZ90qeW
Xqw+fkWWkPSmO0iByZzVJtHYVkLA3GAuww+rShY1ZeiWFXdZT6BQxWJv1Wfwp6olGQk2RUFzIXI4
INeax7wO55tLh9xjgvQfYnBQVkGZ6NUS+nCNEuTogl9RS9cn2J48SxYFGkR4YLTH7WdYQ8GJYi3n
W8BKVaeeY96RMOJZmcCWzLiwBG0psPYtMWj73Q2dZ4vH8zb+vcRcRwDvODYE/NHPdY7W2+hq5wFW
UTCzGMpwyjXt1B2YqDptNmKAKWtscAHiv0/KP/fomJGPd8qzuRMY+PndWIl/7wPNGPUrzEDZn+nr
VmR7uFCQ8Qb9KPuBs+++C5ieV5j6q0x+66lYf8qEnoOOAma6cqQdGB+1i1F6VZbFleBErMs727ku
MWNHkd5RRCDhP1UQgKxf1s7itGlPFB/lZTV4tFoqbI82xSmQAbbFwOCyz/EPgYRKgi8QCq8hirl6
Z+vMviRvuw5VshVc5hnkuj9mXIXmVia2TiuzDgE0RKp3uHpvyN9Ajrc+BmhTwxXBdMGK4hatSEWe
UE/EYaencHcn0dv0f59lC1ICGjxq7Ny61g34Nu1S1W0+scafwgLihgl7jH0d79vlGoeM4nKqWUTp
fJRnRzyAYAWmevBJRyLwkUkYh3blSf4yKGEts3GiIBWM++uWcAEPvyAUTXBuwiLjNy3nuk3ApO+N
/QubmCuisDgWOhRIRyFiefJdWjmLKCZxCQjbWaS5H5s+jJOCiaIGfwo+eQ+DsShHeMZ8kMYTOfJi
ldNzmUNPfSEEm/TrWGS4cMuCw18V5mJJwuOUKutCL97LB0cfNYYAAYtG5GM90DuenGYbnzwkrvBy
7VTEC00hUxNgP+UZ6qa5/9UEsbGvWDDEV7ElvxufpRvLHThscZxkpBO+NzK94hGFE1VSsuhzU+jg
5NuVh2bIYW3VByuLsS+eHJ28IzfoKfjKk79Lof0JUh8h00Ze9RRw+cEosQMKmALG1lQzt7Io5fMr
2cv3sxu6Gh/kIUvHhSrLr0Ye7Bh8Y0I5urgiieWF0oCVDMcEM1wPdkJTJ41sDpnDIS+RVg+YS/Cz
qG5t64pu7FlP6+mYgvv+AZTW7ZNmS2Qf8hergPWa/Mq1IujtKZzxzawWdQx7Ns7+6dOXJZjv/uWj
UPJJUZ66OYiZfsxbvIRIgVpWS7dG+F36J67cZdfZaUF/3g1iTXHi5wWLCWYh7zPRKEdnqBUqfnpm
GzAFOD7R48nOjAUoNVm409cYGFd8Sm4sfnwveKpWw3UJviXPtOhf+BOtsYebUnlL5j5fhx5TMeqs
355Rdii5o72SOWQzbwakgOKX6vDLalAKnNLiP/iAbX2360pa2YTQ7Ue3KcIs0Nzu8ezz5UIx+c0j
D7BiYo3FFYIahK9DzEK0J4o99tebzHpQDZeFLS367TNHKe0MhEeQstT2VYxGqPtrNpbg3+ECI8oc
lsWq2OFgHn89aNnkfQayrrd1lQneHMtr+NNPqwyQFtEKlcrdkJGm4EpR3kPZrLqEujxxUMso1NA6
NmVNU0ICm6doenXh7ZwnzxdmgkqLi9FBAxCkSq6dHPVH3Ve9D+4+gSz9frX3qwuK/B3KQ/ra9I9l
mhSAl7dsLI+0mCdHzXzSywugtH9qq3SFQ4sgx/0P2iYnhtfg27Ew3ei0tsmJW52CTZHHa6fTbbuW
f/juok8RL5DwR8VP5RxaLzUiI2UDZUjzJPObatM1pF4QqWNo7/bckMVb4uNRSFfQkzHgm9Udw6FT
IG6Y54ooVVcE3jSnPx6m2jm+3Xk0wDDoYeUWXe5ATt7EaNcknlxi+xxGCuq15Hx+bx+zmEe3ixI6
dniKYIpnTBbUOPx1eEzDSP+i1EpjcHn25Y00nyTWuh21BI40+HD5W28ZcB/aGZ/9q+pFndgqmMad
qZOlSdoLPbF1InKmVwyYnDG2m0DWFjTTu8m08YuLo1kfFKqN/ZsW0+TQqkU71zBmIHqudJIWP+ob
ftWNTk1k2yiPMScvPU4f6WAabujw5pwY8NKGiT2IEKwelIsEDefLEU2LJ5K6cKgzKUwFqk/fvgFI
jxZOqKtASbK/t/6kndXHjbsso/qxqQec5zEVUYYDqzR+IO3f7y0KwgYIkxmWBSIzOZ7iXgMNwTGm
Y2rR7J+eK+ZB8UWvM7uGbVhTo353SekrD6UugiISRx2QPFMOz6cqqFyWLG2IZojPsazulShEO4bB
075AzQK2CHs8IEVjoqSGLea92CNgiR0zjKvb459x4gUzcZdboV+tTufnc8gfKT5RHLHZmYfCkwsp
ACgrh2m+MEchDsgSE7HPYFr3TI0pmXRzzViB1NTJOh5X5oXjvAYcPylboBXHttC11TTS3w/Bje10
hRnW09FoN5Qg/z7jVGNmBKHF+HLj7FML0P0AS9DUGFqdRrspoy76pVlOcqtXpJYUWoLivkqmfecr
ZpKZ5bQHI89opuHAFzvqqcAa6I1jbxYAFgc9lPyOQPBzKsnwTZtuOPfT0afL95kW0qNQ0109wYau
LIuzGDUC/sJWNvjD5jNHzOKKhf5iNNkgy4i4PjCrFSXf30c0NMak0azOzEAb4HrOkY46+ssOxgLt
I59Ml5BRQlPwz0Ypjmw3+x9U97q8xfLo1nkOaL8Xg7r8zdojDc5g3PjH+hz7bW2LDUXMWvmDDvqi
bdtR/elU2fKNo58wH6BjO87pLsMUnuFRYE6ps+kGxjGowWWchATPSJvcsNb9nBGGfrLZ3dScs9qJ
nljBBZC/uwtoPsCp6tG/MzEvU0pWnMbjWE0eqPoeooIPNVtweqy4Qr8N67rUVFMUen+4Zrv1niGR
9sOk3BEDM+CvYlHVoT1xlvXzVlaR7lEA1cZpTPBrxhyMtaWVXbAMcha55kgugUNlIS3I9d6FedYr
C6eCjIbYkD6NDxR0rMX5KTI/8PD8CyvxnrfCsZN+0fc9qPPZXR86nEMkMPwVYsH8j0HbDYVRYvNF
GTxhPcOKPHvck0d+6KevXAgroQ/3hoK4VFBK2JK9yjvUjAMOpPKJ+6+zrms8ZVzzWtHbsEmcbb78
L81k+tpFO+rVm8XhD1Fpvrsyp7RVAELUkwygX9HPRwLmCtNdVFcW28+M8ubwkxKCYbvv1lgwPwn3
UoiCwjx6Gyf/SaRdetxswnbNXrGS+i9cl0Jbbq3/DGM3Tlr2Be/xO9VuRZWFbt/ny8CC4yvu3SFf
d916bPLECkumIZpzmQCQ8BlH/Ti65A1gY4lox2Nc9MSxoYTwtiCgU123IrtP4jbgehmRD5YV8jp9
RqU1in/t7vVnJWGBBTSkXL+drfDEDqt9O1cXQyR6PBcRov5UAP9ZGMPdTKsZ3+MOaUggJFAVKx0K
mVQZTtkywfYHyz65a0LSWx7bZG9CuxvJBW+0arSqKQWN2yCkb/l/vLD2lFh8ejIFthxFg2tYOWpC
HrL5LX3elEesZP0nNiaCIS1fIFgop3sZuBjGCcLMOOTleeYmBE5u1HzBBYI0ayHvS7nrrbJdNBnh
YEb+KMg+IdF6TBEhyZV58rd5HnneyWbEw8HTRo76IAMvQLhUeOX+Nv3sNxNrujCbauJp3E2xc1pr
cbDW6RsFGMaWTjoXErwFWFA8hUrDhNGtA35j/Iggvg5M5lTf5TpqA2NSmR+R/v/o8sw3ZYaYxsUo
M1Ety+ld8rMr8R1YsZNQOup3UhoalSqIiGMnZPH93xIITIkG6lFILeSHezUP2IYYkfxC/ZMvhDyE
CeFApjjBH8FrxqsMDwsyGuaU4ATe9EQmEE9n6u3uTEWeoN/3flwLmWGNpqNY/ZHhg1PY8BvAXhuf
/uB9dwwrU8v3yjQAMlKIBu+jzbwSBi5pCsbKKiGIOJT/q9cLozVZTraKVzYAcdwaccSbItz2VRAv
HViGbaWwUB/nbiIsUCuEFpDzFyVP8HQA/padhiiFnbyp/t4sea44Hmj+TYo4gzclnPn3cHn4GFrf
YATRK12qcxA1kCVoYypNMOzj7f9zOV3MwGCwq9ux0vO46MHFoiM9fuuIUNiGoYS2xUTnlXa2mEZA
0R6qGCP+dDhosOwG1yFB4fYe7u1oyTp9yOF5VLl5vr5cqpn1ve/lFkMOknbnRx2cYY2mTG+7mbcA
SdpqKz4iLRJ2TX5ucKf2PkgB3Pl0t7mgw7XmlTxsUOB3ti5PR1BhpAxWk4Vtp7p9scwDNwUTMJAv
Uayh7ggeWrhtDT3rzQp6XTstuw3AeCk/YmRQhL2PmfkUDw6HS4CWJtCaTImSWdr2tCqYXzVDzdb7
4CRJWBx0lu2ids5T60KlrjpNwZtNXBkkn8u0XXOLCemh9MEaTCetHI+lVz2Kv3keX7mxjeepXtIh
yWSjqouuiXvyJxWKNo15lY+le7Z8Pyo9y9B5lQ6Kytp/L6NhAYAyzRthUJhWZaUBiVOYjYadb31l
ntFZmcv4J7vIedspKQL9feL2oEzZeTwVSPFGinQJt+4MWFg5MwGFFORiwHD8H2pbiac9WoCr564l
1teBJ0SOdG7Yn39kPj8uj0jD8fI5CuBdr9wEynri1iNqdwkbYudLm0tguJbTJNt0VxW2DQOde9WB
VYXymuV49Tv3kKiy5yrKcKy/n/9wlcxOInxbOCIXUKg7LTeZA6bgRxHyCWjc9j+H7BoVDte+JqFs
wXjSFMn9nhmKIjUZpC6e1pecK0jnH4XkvLYqu+KSvBo5Lo+1hB6qRdAyfTxgpwMzPl13eq2UaBpo
60od4QpH0ZbGfWHB/7bjm6EJkxaxbdMQdI9oZiwI3kSjnvYLZE3cQ4i2TExXbKdc/S4WN+Hcw72O
IJ7afv4uYCBbipOaf7xaIpaMnxj8w76UVgXOgjH/X45iEh7HBBgBwgKDb/cMcYJQ9JIvcw5nc73O
oF43Y4/LGBJsv5wFjjcieXomGYof2cX6eLOGmztJUq7O811khhn8BRoJeLkcC9YJOs1aliBpqVoi
ZyyHuzmT5mQGn2FZKKKXjzNCStf7Fo/HXVW6dty2DC58VRACPa4aCAiijtJQ1yyF/f684t582LHb
jZdioi/UNQ+urxovVPfZWqowXwkIMRn1rk6rIwjJ+1vEcpDCQVvZ0WZRDpeiRwJ/Mj+5YPxT9sZZ
+7akZ7jmaDlZAOGRLFEtNdhCL1X5cz8+EcKL+RTDl9mct0RyvFUdmddg3hlanvb22nNrMpA2aVs3
3eJDZhzJjjtmuiDLTCwzNHOf/eu4ATI6SbLia1NB8wPWe8rdQxtBsv5XHx/BLr2/VE+ZGPsQm1b3
k/NrUjB5H0kZVBQWo9GOtFYaMePdp8/3Tkamef5dzFd+U2YQ6QEUKfRHxfJuWjrCYZV4up54wWzz
4zsiB9W2TLwTdle/vaZbuILhxK3wXCLfvlPV+NTe/Az15Eiyx19mgbR3P0J0RdIZFQVt7BcM6pa8
ao/Fv/1UC50dvelb+MAQuyqqseeeOAY6UmROg5urVrAJ4fMHwRc3S0sBf4ZjrmVyghgl61NXO9cT
4f2aBjpEb8gxfOCYl1Qhy92IFy9I4waNoDHF6XTGdXDalmEffDoGwY9fYfjusedJG9y9Z5lCNle5
ZnCl7gs1eyGA+DMyIJ9lX6KvP34x2/n5WKTfvNSYAR6NinoJgD8vxlSblS/nDbJyL42u5nP10AU1
Cq5/XUgeQMAsglORfQNRthQQ/jNQ8KfvrgwFzdpZU57j6hVzz5aBSH1OXYjrk/r6mC7I4HsMcoeS
qdQso9H+jAynkufsg/5hOTw4Eksu/0B4AvNVuJBQ137dU9kXw9OXC+4k6eglks1Me5aO3tSxQtsM
KXNG99HQsejQ2+HSi6h0Ja/OOqR2DatU1+9qyTjzp0D9lf8r+F1J5YHZ/6dN4JzfF+lVXVbmz6Di
Rg7UULvKkfze/hpgNRNJvMym4Whrzesuw4syzttH/RvQKw9S9Dx6oP8vvQQ8j9QtvjLFZ6HpkRsB
PzKQFAezTCUV0L4xbJ1ImeLNej0tYLbdgPe2z2MsJKyVYeIBiAj/Hu3YhLy8BPyCSWX5JZ4IaiDB
6i75jn5C7mM+dZKP4DTLIpdczyEcrYanzqtwbiDtcml90XkgVAx2WiAaz3bhDNqlRuwpS0v3e88R
hmocGjRA3zH9zn1x9Vr4ecu2ms/0lUP8A2veCUGmiECoetOWVpoPvg8DLXAekee8ZO0WvCVhZdBH
/h9Y4egMiXpuYzJx1Id6mSYQ2DC4ZxkS4oV7/p3FBhItRGLWoeyAm7XMct4Lg1o2mIwYa2TxxzWo
uMkBKFdhC1P++eAaFOmXRCPr3C0wmrCF8H2MRl+x3Y6Bwrcf5VoQNM9CCAlAeO9GAn0egA5zYtAp
GFyndL1vj7R+TGlyNi20x+Ic8p4IPLRFtiE3obgYzbmK8n3mi6QTjCRnByqpQH08CyAuHs9XtgW3
WQbu5rNq7gcN8f5kxkG30sWScxNYpL0MqrT2zFSYvDlNz4iEVJalbTiJgbNEQnm6rj7/wYCkiLJu
5i68DedrOkM8GzjwBH/nGpB61Lg5QZiqfqv6Euos58UAWbTSTiDvXLVB92jgPkt7HuVuThTLXY2D
poI/VIvI1n490I382FJGq2ALYf1jwuIO6NGzaPP9rAZxYFx0teIStlMjZIUDSC9VtA1b0v3G9Gs+
0xfofwSwix+naeOS32Voaj8yU2PdHdZItgvtQr2el1lwOMG35mjNNTvwTyKmCI9oHFrIaYaN+IDx
1vUEp/dOVvbgFJlHaYyXK3WntHcsdS3/SqwfQXnQddU1tuB7Go88zIhdeK+qIVdFtMwLrh02+1RF
WsNOfQvBXomsQdGQR0N7wSNevbiA72dWr+6oyO55dn4oxURUdDTyrnZhKsuJ2t+MB8iQd2lRksnW
XlbyYlaWiojil+XUJ6DV4dB8iExdXtwz3rOB8TKYodxMKvjw9F6Ji1r2TqP1jbbZ1yH6b16NpixL
y59QOXhx++QF/SHaE8leGuAts/pYwbwHNPK372UUg9gG7RfwL54Pyacar4XsgtfuI9v44nz56sAn
M1tVaFYcrg3bOxTjRj+wLiVIG9jBlGa1466wlMDx2PC+xHa6A+0iy9tyz9LmMinj0bmswl3I5PhM
szpec9GKWzFWh/dHDowdxK6ERLJggSepC0RbwvI3mIdHPGNAK5CDCEBcjLUxEzYONuPKMUJ5JjSk
M1TDHZqdwdDS7DNXFVzhNxlfzwvGOQDoNg3bTQFnpBvTkFmbqWo6tpyIv25iRfV5RwJtN4GrueAU
XvPJrK1tO1W8Ym9O2o8rAYfGUaXmUGxK8vg23jL8euqJyVh1nVzR0s5OqBAUMgF9qZMnAGpWtKzK
SBCY88+YuGP1Gh+2XHEzpd5L1o8l2mjptXv2p688vmZxW8xqluXLnnitfs7P27sc0Ud1efspH1xF
FLYF5qv2DcKYUqNhbJCzl161jEKCu5p42saItW+GFnjkC0FuYXRv+MGZRklSaA61Aan277p2S+W8
tUG2yhM7ORnd5dV6PRS34JqrP1KPsfw6Qw+S3ejNX6pUGwtN7E3aVKUfJRpc9d44N9npXcACTfiw
Di0zupDeVtKcB1Rrkf+sgghzM06GfAEW0lFCjTIWT4cYX/DmUdzgoGphW8O5HT+9/8xfT8x1iqIb
ewnPUgYoUr7c7/yN2VLogNfIFiia/WXfneDEvNmo0UXdQKBh9eWngpaHKlbQot6DrTuaPLNpkCIf
Xmwd0KucQzhgIv4mkS5OL9KgX+Vth0Gmr9rORRbuv+MvMV7ASZ97GCuAOHEQs22Y5FOVSx3CdAo9
kzolnVmU74TKgf3PyilETGorfIOz/k4HC+eFcQosdqPhKkOys3KvM+AowzFKy5VFwNkmN3goah71
cqlzuLn1R/eNnAEUtsQPQInyv9kSRvNmg6RAyFuYtRsy0imt903H64NUdZnVKTZ7EFwMKi5cqLdi
RGtyf2MU4aMkqBqf1ArznpZBTFA5rRgCEbodxL67z1FOwq43v4tn41R8pJor5knKlVFn7nlP2zPs
aYaLElWgqLhVOPkwKmfzPTT+Oi+072sagSzb3VO43zGLfp4Jds1pFY1hhfE+eRT1rZbgNavbtegm
uMkr4z9Iw8DnYVjPHjEF7ZA2J6e36LmrbgwPx8vwsa9ZXVuOKCmrrqVc51UDtUNNepacYP/83nZJ
JYlBI/hHN0SXXbcutCz9sP2iwmfVyPeEEHY67aC8P8aYDriYuO5Y5pnNUJWZDP6+T7zjTNl7aqEu
1o1W0lzX1EtYkyf5upM46LX79SpzYsOhXqc7pZUWC+YUI0tTdNson+s9NRDlPcK9nEKLx78gE9EZ
ZXtBBHaaNvW/JGzGtWdwChg84H/hOpRAqD8DR0Lxv3e1obyGouls0mxXlCT+vO4FjTtdbMtCikfL
slO22In/87zHRK0WC3ptDeqOC2Y5RuTdTdq+DDpkmo0XHrofj233ByhEvXIg0wBXeKhlFwonXqqG
lvKdxox2QAT6VsfLVXHa6FQx8hqNUibl3LV1wDUPyt0XliCdxVfJ49tLVNBhQzhVcMyiFAXj+fVe
GJlgiHotnftt8nqejyOo4bNxYCVnnU/WRUMgvg/0IXKBXYGVmqk6EDA5fzJMsmhJSChsoruRwnvB
QWGU9bl/DObRagKruOY5SoAVb3wXxb0gdGIvSvZj5gI8sD47EYyz3T81bnNnjg7j0CGbrZVZSqNN
vS+feqbkz/8MFmD4qHeEQ6RUfODRnUh2MHbXBxc3WE49QmOKepqAuLBhtn/OvwUaPjVNwNY4jaCY
wufniBxS6+HOpci0kppNYuhFSwolqImh4hYcr+GlYgDVuO6866ZfQnUX9eNgoCKhkopcSlHElRcz
GWUwTcxZQRCJK6vl9HYkjycAx//uUvjFX5mNUO+ZwzYkMKAAh7WGWTdVnF45BWrsw1ee52Q1C2Jj
UbhCSjEQGnkDjfmxeVvJBpRhk7dMaJl5fC3/mF4jv/zFIkHhdp2Urf3SVZkdviWZIOMTF3fhJKFu
8y8pOgORwEpAEiHknp/Q9YHwd8SJEzPwXoVIV85GxpJrgg7nHXP0sGOqnO7EdWSIDVNWgjo15Yv5
QRiW6egV5h81f8BDowEeM/zogi1CjTVxn6qKxlfqYPk46OqaUVcTv7v3xXmGT8MUJ3lzsFF7X3hN
Cc/v+q7q0Mx+F/0Gqju3vCyKJxBN5qolcHxBoz2+K2cva7vsxAGy8OTIifWSLzB96wYU/qg3cGV1
Jzj1EZmB4XWeNmK1/phhGfjPNN7xnO7Zt5Ef95pcPBsKa5WPjDxgwmFOms/Q5svw4uVqFdTt7lC3
7Q4HoGyqGxc5SpRPUXwws58uk++dP3RrT61db63vnCbTH25mhjHHsHN74SutfhetpTkb/NZZgazC
LVJaTvG3LXZPTp9yQRCqwtzmKuiVDzmTf7OLoZc1+YZApledurBv0Q5J//dgLE4TxC8BBLM3Rb4f
8b5aJNRjsy3+kP1atn3olXYNGBPUsoXsmhIGJ1mnPmIW8qG8/r3/QbiKQHQQGK9Wjkq8IxiVrhcr
cPZSAMTvdWG/bh2s6x90whgylcoaMSlygQ+Zo9OsP/SqBw7Bg9LjcdhJLJxTh8FAQ7EyMu6ZucdJ
3FxixSE15N9pVb1XNPueGwa3OYIRGtB3YKDnwPjV3gyrgVibltZYU0vimUQmQUOLHwBmGswZePVN
DvpipCPkoOnE615+ml3XRsdQLS8jhad5lVa/4A/WKJ7riQNqyG+nUPEBSQQTMoffpxoAkcQxvAqC
L1c06AQKL6l9T6pKJx4XaI47xnJUMFKyjqxHxLVHjsj4L+YH4Y3f9GL9piuuAKO5cFR81mC3i2P4
q6klYsFkrscMSTCG+3TghGR9rk0yuUiAHQx5WKLdLxNINumeACoZoijBOgWiPAzP713Lhdm3LYDr
hYcx1TLg2YKXBdUXjL17/IRYxId8ktDFmYwGSmXXOlerNfbg++tfvKk2Nt7RO2uPgIoKwdkox/LC
z0h0O6HEO7c6ADbBO6Bmvhh3uXvk2ybRt8IBY2usLc1rUdABRGI6M3Kmeq8FtLnCIi/qrZbIGhwn
SwVF8fjfrm6pg8t55T4wqiufgJp71fuDtgzuviHVm9xPA9jEvD14KdNkYmzbvVkKDRdCmw6RYLXY
Nbb6pwjk0hyn9Wx8CMyI4cgHV+g1i3fZs2XIDiQbThPV4UMi52Ed1C1oo7KbJZy3rK6/i2nBL1Zy
l4fyLlsuq0rUji3cU+eFSNF9xTy2z32Sz2tKV+tEUd7yQnZFrelHs277atxNv3Sybr9MP5SIla5x
90Lytamb9Fk40DrLriJoxbAYkOAi2BEA2Td6H+Hg6pTF8+3hxWpUEMnufUcqmT9DGUCMzhTB9ujq
J+wd76HeC9IvlOcUUlRcTUWVUe4OHA3ieScs9of7gQ1m1m+Tf0e/Ra4cJQd5gxrF2zBqdYj/Nayi
j4IDr6gNGkedapC25y3/307qUuGh8/6rrFHpY89b0j0LZQMhzkpO7KcowgLgvKc1KbnDg2dk/h5n
fuofuGCT2oh7PioITlnI2aNxa7yIk7Os/Kf59hgZVbGEYY4LO022BQUTGHfEWn99cw9zveOWcvXV
1jYwt+9QvHQhmlSYv73DHzg+a7kOO19V/VwHSmrQ9F6twEnbllN8h2Frg6Hz8mfYbAuARGFB5oRs
l1pp/M2nrYx0qGzerejC0Pby2eCh05vUkAH9DsdPFTpTvbccbUX+krNYRAo7rxXQOtG/afxvsCBi
4XGTSeG7AqDgL85UEpy+pv67NjsJlOeQyUJdxp/b4Tbay4A9XnVowtdqfOxEmSA2Qd/JYOCVgW44
e2dbJlrvz9jy+g/Yv7up4KSqOyhG+tABMKjQL+UDs/cJJPwpNtsZC1QH15jzbKaL7iRurY3LTRvi
ZIQpSNovRcZ2vdWfPhruICwfW/I7m2Kv3eMihVEXOi06NhO3iKXulZCgLp/bmmuE+p4PynorRVVb
qrN0+bYy9NkwkL5owRB1xJTBj2S8GyqSlhqkMdEkFhiJBz8dkGTat735jVUmLh0qDdXmkyQSIRZD
UN50U6PkJ7wDM6fSNH8yAqsIeEu6PI/0wlFf2G3kG0E/ap/Tgip67iYI0JjjcK9i5YBSVUHEmVjR
DvDyI9lPJvJp9/srGICY9SOFgaakl7D8gIEbTI0ZXVAP5+Wj84KaNfImWmeC9wKZ4x/atnEd9C0X
X7sDrCPmlokt7/4Yt8wsPBYCBgm1i4+vxcXXDJ0MIw+50iCQzNRkyMVuq3mSfvNZT3hbq7H00VE/
mOfukOgpfSV9Y75ZV9Th0Cx9o+wwHjy0OyqM2yl9TZjyBrwVRvitxQ1L750Zw1prPgJRiDIzZzdP
3azPUMPswe3ncNWd5T/xBRCFNMVKwNaWQ6JRDkr22mTrcjfoU8tzbe7SDzLTGPwtUn8DX08ypT+m
YFEksoE1JlwKOJR3m/Akun3K8LRyYBQz8BwQ2dy+yXhqRFojYy4lb4Cqnk3cpx8l6K5fJFx1V6Ip
7qqwr7MfZLvqsGNo+Cu/7UHykBpai/LJOBYZ+yNf836kmURtdlAo8O4eGX16etLcuqWIqrLwcl9u
0yhfgpMUZb494fYCZVtUZ9sJeFfrny5IJnC+MKoxb5vT1GdfIdc2IkfWgwld5Yt3xYpYfrI+yhsJ
Kpmw1Ju4WMnKIU8nbuMy4HBq9UILeP6ghxEjKx5kwIaFjE09ylkQ5nvNeKXHM+/LBYaFu2XpcJbA
PURUSjmVJutqbkqrnHsJGnFFbvK4sHLpaRITWuL02USiYKQhNdiRDppDj0xdaavRFYiEPJvLfnfR
cAg0nbl9nxq4dV5y+9DWYH3hxrMYigbHZoWHYjoHNCoEmT+62P8tcfiydSpdrCXjxwDrSiBhWax+
sXsdMnQyWTzP9nU+zSV0pD6lYVwJEtKVTPtPLBQ9/ktFfF95vtppzVzxQi24YsnrsPmGa0mvnH+M
/UMDjQXWANfq7mnuPjUoIz73BSJJuD8AxTYva9Y8n2ZZWQG3Dlq5Mp27K1p+gxPiEG0tPQUdrbyi
7iW03fm5vzyG7w+jIMDTSDggr3InaLXhr3e977wYJGeyXJDoc/F47fY+s7SL3Qg3yGGKTU5jU7/7
Gmr3KiduzqbwtOkVw955HVfWjPsOfMTQm5txJs1kdak06ULG7fw4E8kcBqvfU5Yf00H1gFbwg6by
IkjCake4oYJSw/T1aoIN7P3PX+AuaCFnyZCr5Mi+wk+Av/Ka9v00TrgKn/Elgyn7JdlifQhFhF4z
bchKo3rsN+616HAwaoCtTD3xziabB67qbDcv5rCql9hA1s9zJ3V8mNbw7Emo4SdqeVtbb19Q+D7b
F4Id6bw7s72sB8kmWuyNmq3P7xdtW9Gb87485rWLoLGfSxEpJskOHbdNGtQ1lEiXgcWTk8/g+ZBH
s+kKBvhWsJAUZV6G+6FA+bkjkP4WUsR0cPdNOiAI61gjEmm3oOmkgJ2dj9f5GIQ/riqREU+zoFNE
X1HI1sByWFucVs/YCP/6+D5XY5tXo1Aq2AokZdJjfc2Q2yaWAMgFbmsBl0Mq+d7xkK7TBB3e5+L7
iyK8QcCDBlxYxkSAEnN/tyMiUaF/QhjWXwLCYnzq23xBdOMKXT5EDH7hhsRmQnH9GcpKDu7IMPue
/tHTYRnkTvuDFRMg5sOCOScshUpAt3suC8gYTiuW7anj/Tt/jWgjnbTAnSCOPpyC0ZU1zkZFG2nc
mS3v1TJhnu782/dAPl3GRDjak62cMVU6H0YaqxhUJ8+XUpwbW3ZIv9Ra2U4m69AE2/NmrEsz3PNW
FL9pgiMUyLBRROLDr5/ppkuSPflRcMJf0Z7kmID7SnKjbL/pSdtNGXpIrP7qqqSau1KWDSXAR1pq
LeCBX4WdlB4/6tu63uHvgwLYOE7k9UE3PpBWlWrevcKCrZZH0kr7R0akEXG00ORaPW0pjrfntkgg
qHgPyKFoGNGpdDBB+LlDGsRs6ZgBuueZFUa+E8hCXKF6aP6xRHMRsBolOntuWxnposTBkKUlRQzA
fvbfJf8mGyEfTv7SPpI9Cruj8iis+02eFYr88dwYH0ATunZo7Fp66WHJdpzSH3yenOxTNhK82LN3
3+ER5PmSl0c+Faj3dHkk+bdYiSz+ZM8QUYT/tuyKhABUIS9IYLmzj9Op9E3nDW8NS9pEeqc0oO/a
eAgPdO4rBIh4n3N4uzGNKnrShbyd1kpbPEPVPzMX0m4AE3S4OzC+fVW+trkqqD2ucvhVSVLrw3ed
n/9a5qyO3AIBq0LNggQuhbKxs1P7sGAkOhdBP/A/CoXXskQ+GBdxz3sz5cC0AwCyKWoc6NrFu5Ft
VbwoqN/67EQ0GR/BYvHtort2EWhb20AHormjhRWEBeAUcuYQ3NxA+9IcT4ReI26stFKeOwJHp9Fb
CnZXt8OQgFPCrXLtlZqFFekHoTOhOCXw5CLGJjDHuz9MzCEqc64sI9Gnbtmd2rhOVAuAYdy0zs9c
mzuUCL1QABpd3Wm2DRixjMOXB8TzK9h33UaI0ieumc/d5RdIh6CI9kTcnoeqe9B5pLQzO7NIogwg
5i17ZTDkaAYjmv5XwdsVx2oomhGswAriD3RUQfdwkjjNKvVVEckc3HC0zwBWQggkRPSEkv+T2dFe
uKjaKmwTYy6UyEUxwupLt82tT3eeYiSL3BiCBFWMe15YiS99epzGpnCnDshJ8pgUn+iyzPvFkTQL
nFCj0/WW2uoK8TG/blKXspqyVcMt0gT+yILJAFoV8jW+mfy9u4sRJHf+Ht9WA8WoTGoRgf1HN5JN
PFhDAykPvGjcXtYlQ+XCeSWg9FR0JcEWd0SKPe3of4zR/Es3xeM8dfoOCx1KXi2PBGCRAPkQw9Wr
Iztr7uNip18HvhhE+8jFVu2OlGIIxQ/TX0h86yiDuDdu4f/i2ilO8Qp7iRWSZYmLBfz5sqdw9v76
ddJ4ERtw90uK0Pl4lQ+OsXQN8DIvS6TVEpvL8j3OJ0ZK/NS2P5o785zCegiIyGP7/B91Jp3Ty6qx
g6bf2nE2cEXu40lSrCBOG2LqH8pk2tcrK9V74Au4vD0KR03Y+gkrzX6L5ebFQE9n00QvhX8jfaY+
HpigOJ1abeSsaI/dgklglez+UTSDkadbQZ9yeCkOrlsm3gqJiIu0fQCerQwIwlJiFouMJDCn52Pg
+Jj5xmFfNeuMSbXKPtlEVsRqZpOZLFBE+wBYNGXCm9Y/zcJmTqI+S5beD4xjuqWZaeEP3MWbuIp0
z0CrFOTDZur+gcVjX2+tAtad/sWyDSyszDUYuuRJ50RVj+mvZJ2kNW9nE35ksdP6XAZUEYORT38w
9z15LarwJHwzouR/KEBVtmdt+Cf8LaUSzonIAnCavh7jKz5T3TU73EiBxJDqHyRTVgGCQZ1DItXI
qV0DY7QNaBS4794uZLuqQfFf7QmVvSM+oBXH1qhI8V0iiToz4wWoerTbW+flYZ3cqdtocuo+FadU
Hk7g7koPDl6vHdJwSTGHiF2D5JKS2huZNhn6DJbzZowk6OsrB/6nGI+CDO6cqKGgiEJS9MAhX4/U
QSR8asYC1L6xk4ZoPUWyBnqdSslhulNtwp2cOhr6aAWeKLEvj998SXuajLJY9Fs/cEnbonsMz9NJ
JeyzqeEQHkeG82+I8BGtnUDu2y4vTJY0sQEuMeipggRMUZsW0/eqBE1Fm/RqP2X5zdOGBvUfmLVA
67zF71BS8VsO/UKq1iqjP7qRkqrK3qsA81xOJEF3qrCe43O+cbVCAVuxog9tEbr113+92K139Ekl
kK9lofXnH97JXjerUU7p6b1cubMkMqEpOboPYLYduVI28uoZ6Xoc+Ux3XDHkH9HROmjXL9IOqsE2
DEaLk6Bp+M7CGurixxNNScb+OnZH4Fq2PZEbRsGjGRRJz/l+N+T/KckFx5WE0ai8+owv8STUtoxH
uUpMCaxljeIGirDm4wphJCQMv8yXK4EsS0p0WJ0nKeXkRgNVt1rMvZD/lGUqxI9h3rQEHksT2Q1C
j1sVeJG24fNM+rdZW7SToSnNQtGZ6txhtwuhJLD4RaRzrjRuv33Jrl/Va8drJZId7/2mp/SqgglA
EcCabHyi4wTyAGnK39MBXbbrBtwALcq84BgIU1rHZDkHc0XOjXh2fQBpV+j9mqdOsAjk3Nklq+MJ
h2MI6nwqyxYG3gBdBNu/e3VIFleoU1uKc9Oma0L1ZUb20rVCUSqp0+ym+lD1Q14c0vRnc4i+gk8W
/z3xD1m7E5vOyc/bqii/eiWdJeu1Pq+OFG6IDA7q2aY8kDUUJY5KiFn4dQhobfKJLvhZo3OjohAF
pf09O3qW9NbcCnNdxmtoxXCQU+GuBKjIKrE/7aCmC6KjXFfXkYiC+5/xEdYvLsm9dIjK6goDuLuB
JCyb2vVaVlPY7tywv20vJL4l7s6sg1Luhk2aFVkOZDqHs0IE6smlhZJdV+TVP0YgHTLbN27SY9fn
bKQzkNgGaOkQLGZDBVQ/c09nazepo1gRmFTc8rCRyD3KzAtBt3ldmTHHeBuSLuR8BdsyM7k+WKgK
WdB3/hvESIEEl/IMqBvTzJxXo77nHn46qn4JA/LiFhxZwE0gjJnGm8tasHEVgEyV9rVn+FsZpzDj
vf042oKrV/IUl6UCpYG6LesXmxUAZOrHpAY69tgWK1uNEPaz2aaNoyIUbz4tAHUzbCFF0iWdhVV9
7pNlCSLjKCJRdSykdczQPbPA5rQfJ0rlzdO3qnYjn7DQSKOYcm6lU0zxAYOINHlOgXwiQUOGSa4T
RtOuy+ymrlWyhV8Z/xsdb9iOJRIeX9WUK6s9IjrpjKyF369lRP8ErTolLRnEwKrk28fSxbg6m+Ob
bKS8me0RQaNPmwpAiFqVbZSTCV3lrXifqcZKlOJuQyTARXi74/B28ER+1EwKhcrvhPCTILT2lpYJ
lo8UCaps/vr/6gi+rCd6+w+JcSqlR95nhWKsFo+9qPVtoSyPVK8Strh084vU91PbcFapnxFYJ5wo
95Piu8xJR8YYJDc4UiQEjukDnlfb3paLjk46uvN4XxFYLbw4QiU6JM2tDUTYC7vkszE17+x4R43R
65wOaBhExJrp8sk+KKfr/EzjN257/1zx7sR+OdkLT3xKr6XvUmZYuVM1W/rHPT3mrECM6RwonHOw
xTXhsZ0VRFkLctufepW9ZP02IIxBCBsHkcs4LS9FtvwNm8pizSPwa92bIoKOS6uCu67Yi0xmTnyr
FK3DgRo8gJcz06ncx7NFSSD58/VwfCqokYkrdUtdTNsimgXsc+3w9ccom2u3+XR4TlgAvt/3T1tV
rnOrRjcjgSuorIvMI5cWCnfuYcklF2TDFBJiB72VhRry0pDoitp6OTA+CHfGmRPmO0jRg/eAYtWW
NvJ2d32uT7nUHWtNLjMXDEWZzbomI+PQOPl+LZ+fEcsLFiTsOtM4Q5x4VHOhMamM5R+ZQVOY0chH
P677I9iXX+XMph2EGo+Ac+D0/aQX5r/ScEb7PpXXkq8X9Z5eeSGb6dauherKPHyEoYIyfqgQpxez
Jswco4IETrnESaTL00i0yzKzVpDJHIUHM8LWlwUJp4ZjNxaWFKK8QzPNCBtiOIlb6STGmrN8V7M3
4v7vBD7ymvAAY6UJotu+cVGPVXWMITK2Y37IQVxlKW+WvlmZ0Phz02ziz+JnXGBxL/egXr3i849C
ObnqQwNQBWfv23Dz7DvfdAzx1fUAGiLsQh9+VG7zKBsGRc0hg+d0zCBg7Z+JlW+eVDAGIHAAics/
DepuHVPoUFYx5+0oyderzLnXluFswHAJlzHqqjY9LH/ypKOOB8sAt5XnDGBY6K6+JAKDwgYoxP3j
ghwjem/eP0V4lSKSC5Oha2A4NmUzRkS+XZ5izONZfWrv/CIhRVreZv9zc7ZO9gifpnLMI4siYpL4
urbyw8hFQlzQxEXaAajUzw9nAXv1IQy6FkyznGW09cbTT/WOQ6Fnzu2hbvvIXdDjSInVsoaeNATk
4tmcQUZ2eszF9pW7l6miZjDcXkBLFcN8+q818EZdVvUhbw0evI7YyyQdZ2ghfcJAkcTG2YW17dD3
XIqg1fv5FoZ8QPyC1Q6NlSqQteYPPFRbwRsJZGFXS1Fj9F+yzDgWYo6hAqziDQ6OMF77Int+je6U
XBKGgLQ+nTXKj2z7J5zvceoA6YCffcmNlvOWNE/HRQuhuA/X3aTndLobe5ubmN9bPwgS/7L5tSxM
mVClpaXhNze5kFpOClXZkhO41/d3wFPI9lPM//bLXfU1TYdLVTBKxuZgbuuqjZIg/dhy7pg7X5Kr
X6XdTsvpGzzML4GPPEq5tYLOJjeadG+mS4E78D+7WPgQotfwLdLh2E3A/EqAdaRmWxZCfNDqXmUz
z3fMBMMa/xdvD/zaMHoBY6cm2LIBRpKFKE6UWnavgMYV6AI/gBVwIqIBHprPHePetMls3aJXVXsp
98MGL3HBNnKF3oR7RhoIvs/ypjv0FTO8ZwbaBQv0y9lYto72hbbL3DdSKKfQrbVYMUGGOiwf5N2k
yPH8A6QOjxcSUydfgDcJBTCjGNhR1PfaWrBNb5THMFK9rLQNs+v9XI8gnFnttWdnP2kRNlBFS+Nb
3Fbcn6TFNsfipSaqKBz4tL8Uc7YTxxbgurf71Voj5obHhxMjH7hKFRcCZKWgDqwRE4sAo36+e5gk
WIUHjtLZpmvfcZoAstin8/gqotgc3n0FpWuCP6/Gtahj964btFb3x9P4lnTzIQeYORWohEdy2wvd
ljkMQiz2tVxb/GII+68Cp1CCzwPfa8dX8Weiu0rzIZfiTN10q1zdw+qlCeDsdAzv1yk6H2YwDV26
WhWPirCiHvaeTB7+S3gPgDp/aaYInpYdMefGDe1vBcHRweMO3zh/Qr5fgKjIXmUugcPx2z0rmJ7f
4AP5TcQg3UL1ps6UKLsp1Cm2lysNNlHeYTx/l2ARrUSf9T6VCd07sFDcgXylot/1JEk0Ne8sWtrf
o27gDCNgAcDz2wwSEenANYxSbVeet4AHyD0KfaQOzYbCwJH4tmJK8KlPRLJ+7ZuTSa2UZuTW883u
GVfJ7UE6reoXE5AUJ5YNf2dY115Fh92IWeHaA5xqVU3fv3sNant7TyrolaQRChN2CIy7TFdliWWR
dRLHdJ07gq3Fk09x8MRLc65Ef4UxKX9WEyZeny8mRB1f1hJnsKR9MDdRUn05bFoTEd4NgwB1iBti
w6n/draCF1RQvGwNdY50FCV4Q74BkU/55Dp/w38vusWXxY+rAvkUno571R+hBSMPCL98X+3EWZpi
6+XWlS/B3vJQNk9E1u7wKqDMHb3sqGlaBAvxQblAR9DMwSvIMXz+VHgK/HodHCt7bU4bM4lgiKMi
wU1pK93QG+WjoKHGh3pewDywf69rZkmct4DHbtabDvGJ4a8ZJUTQse6UscGHbtuoJxrt8Mw2aUzj
GoxbogOd075lZDbBSApN0VwSvK/dpNKjHe2Ob/7hFrAsv8cxwF8yJqXavzrX9hShngkS0XAsNXBT
O0HiVqWxqNfYaQRx49MtC+bwgcb6LKiHYVCX4DioYfXqb7bY4Wv1qPHUGvNXvvCwW/hVZ8Pjd+D1
78tGkNQ5Rtaq140WSIEgPgoSaIRyrklbgfyvlbMoam2S/TNcAhVUDq2CH7Vkj6bIjeeKgXp/5NjR
2N+vuum9lIKQdgoixBfgLmOqPusxgQEK7mCECDL5xegrZov6msDBWNphIyc9Qf/C92hW8k/QEKJF
Z8vAjBeViMLuJE90bS3PJd/CIL89cmCS+lGEP8WUHlv4oD1V7WZtITM/IY2VDtiVI2M0huQ3s6f6
xcc5DDdFHqincjtPexBH0xlwc7BAl/ifPyn8aSA5uVyS6pr2liHqMAZ40+KALCohtQJP3fvt9Y5K
r/t66T1wu9zTna1pR4QK0lSwvoqx5s/6RzA96GqdwuXc59BdNID8Yl4057kbQ1NBt4mlRhYW6cM5
u0Q+bYEXalJ6NzYZPCTumO58d+gjMGnBkX2B4TXhWs+dpKJc05c1m1lAax8pfqkx/ORzchE1yrW/
TdigPXFE64ZR6hQp9lnzhI11hyre1R7WLyFfkjGshbumjy6xYYtpDb29b0uxw/ZKmJQJZS2aSI3o
x5dianwaR8Isaneq6/MUTfXH/L4rZ7WkL4GjdNpxMD7HIYywBqyTky3w39nOtDKs/ZXRf9EVlg65
T0mGFU9lKqI9VtXvMd0iFPt6LWCXQ5E4wkl3T73oufDM5ilA9jOrZyhRR3ZeFKbVLiLjJA4sbSmV
94jX2Fo/WdqzVpdYRZnyi88puYMhkwn3li/ks7KBuVu5XbejT26MZZcqxX9re1W8ItFL2mCagpYb
3Psguvb8nW/xFZ99lHuDiidEDs9q13M9a1gdnQ5lq96eeNtYdYhTgsfrit/Z5GE254pblkVCKArw
BkZMHH/D+GEUdLM88HW3thT6zY3FjAxgxvDbhUB9IC3ayaJdq2dl6YHaXfVOs38qHQ54UQadS7xW
k/367lEnG9U10p2uWZA7NKmXcOW6TEDosuuASJE9qItBHLMDFLEPY7FY4rckRnDDFMbKctm1rGrZ
JUerRT4M8UU3RBaRfSlpdccn9WyIwK19kUnDW50pinGsVRimyDpAWGBryuzSRaB/vMhYWUAihHe8
bX/ot45Rm+G0S10CR2V+Pq8nm8Y2RV/rzOt/mNYOIW3xJWJROFPcTKSj2T+0e4Wq7cyEjDWZvcia
92Dc3CNw5zl92whDoFTe3eHczvYFJSKmDsV20YsNIxXKP19vLbb7mTBhvg+sIZQIVAAcRGZ3O1j1
hQNNcUGi9Ih0/okPbH07VE9E40NVs77rfgv9p8FpsxdoEaFDmzDdlIfuSVZMgpbtnrTBCLDxgYXY
yTIji/JnI2bNAXseYzAc+ErXmgQJtN6T+Cdnhn3jB38UnYCGigTzwdGh3DNfEWne/johl1vZRZ+s
4SvKm4SdcHAD9i4SFtrmaaI6+m/tLSH3owzylVMnC4UwP0bI9G8u1yfFKPSdZK5Kw/vsdDl8a6bc
WEwGJq4QNO05HBHv/DBSao757NaxJoHTzmqQlPGCr5EWokKsa6lA+yeMN13YR9qnf6CdUPaXSHaH
+6Yie/w7rfkUozsnChuE4IlMtU/R0c6y49TQaQvseMfg0T2vxuQdwf82gMguUWDHl/UKCEEXSo29
ADe3ywggB15h3H5bO1ws8DFXiH9rgAkB0Q1oKieeppOiONo/u8O3CSjaRe9nTlIodocb+Y7Ih8au
bJYt4DVVsbyriExYCEWxa/JyF7hUGOciT504TiAA76b3itFr4ZPoFRIN2zcMZ+NBuBTeFV5ZPZUZ
R0WhIQ+owTgtB73G30NVrHR2Bmz7fvCk9FUiuHLX1TT3iijeHz0e+roAAog0GoLpeXM8qg2vrmLi
9LUqvWYCGsMqfvM9hMYoHBYeI4LXJxuhS6P4nl75rvABQpgCI+RX0Skt/J+ZMmkIdvw0TSXQsmuM
JnvODsDWqLmkVUrMFECasGO7GWiob4aC4XDWSpMfjgK8r8hNehw3rf/qYm3aEAZUMPQ2MgoHBfbu
w5ItEsMMGPMx5okTbAa8uV54hlsc80TLSPxGalLqA1/Rk1wiF5JGAgkpSEwwymT14VeebXz0o6No
4Tdt0EH0A0lKwppIH1MW0sp4D2UTZMKbPvSEJq7mANYrT5+MLPGY6XvjgHloAIny3cRWDenIORj8
M/+aC/uCw6+H93FpuWnS3ItJSKRqZHEfsrKXRJedc/mXYWzVMO3KTs5ARkyQBaheJbAOo9F0uD1L
LAwkg8/TRWhg3sndi40xoV3j6wx/u4wGwc6eEAl3KfWKoEicoA5kgnj2cx21JeH/vIPtivXE9cz0
29tJeCCnFsuaYLdCXszr5wqQupoo09o8AnPIPH0T1n94/vFbtBJ4KI93V7wZvubkjfZH14dh8ss1
yKI8fxaC/CIa4ONxhwaXOEb3DVQOl/n9/XJSveCSs37VITH+fKf6PukocwbtxIy6XMcUQDVB0VRR
IlWDr/vMLE9ATwet/dhPKzjCU4hCZvC1xjjiD//k3QoGd8N94eXGhzjaav2b7wHMuwV7HaI+6ksG
j1WCsq2QOzdi94KMv+U4w8eSZODIgP9y73artVM4TV2jveTqyuRq4dl2SRWrECTh32jnVxh4cwf/
7YfhrjrAX8/UHvcLi+R0t0antl7f7aG0E8mBnw4DKB8+GxW52NLP9oWmlFxreHp1iQo3Gw2t1HgE
C1PQnHt18cCuUn+8BGW0FRnWVw7cYygQ41CFZ0Gjbl6y1E+WjXjnJRUOl9JWpL2dd9ZcPM32GVCS
vTpqWoT3UAaICheonlOtnTjByYICqVnJy0KYt9Ts1YL4K0NUVZYWX3g8BAipjN2l/PGuF078xzPi
xieWm8vaivtATmnv2mxUcbuXVls00fwVK+dRR29DX5hDfmaC44RaZIH6OHfFR+zJa4T1kiqACW2g
xKz3Z+Wau71duSZzVTmCTCMEuyAo5OV/BosCTQ7Uj5r9IQVcCw/rE+QflPQu+pm5a+wilr/c9hOi
t1auphcebHJ4803Wh1sWgurdCdZtLjJyu1o0E4T76h6OIWHtwEm6Y6VlGM/mbv2kdtovW06VgeKq
DMDetwPz0irJtgdjQQYHNLA9WLTbPgd+9UhHI+WuCcBv3ItNBBti3fJT+ynFskw8Hbo3EXyIvfdV
1xOOKV8jvveZurLHtBdGGpX2RHi2Vcb8fBi5pwH20fVjvTQMHGRnKwh+KRFrRCYt0jEcl1fTkyX3
uN9RcjA0mlxHnWPpLBacAdrBISh+Sej9M4XQIeszUzDWiJO/g6D9IQ78/1HgyZF8SXDQWbXJXQFR
il4hDZ/jnofYpMmE4i8/zlONUWtb09tu8C9Nzt/h80Vw20EfwfbgGXOpnyE7RVY2N5fJX53aWGxx
2NpBYV/JqloYfz87ilMS7T9AQdTRkTzfHwdUkwtT+Mpkvd7oEYDomNFqgaLve8Oxf6qzJ3uQqQy0
l0viw62Aep10L/NFFYMYyrq939BH6z7onkk7BiXs2xjePsgWF1/N6p+9ysGBZ5cVmiVSxHUekQuh
lVnh1DYcRWwD5tKgdaBMkgyOehoMO6+sv2D5vgnpxitKhoZWz62mXipbbsM8/6kwCNfec5mX15rw
8vXnsg+utpwu4lZxodKvhMDQgW9Sj4NB2RQp+lf6HRGLKqSt6Z+PPP4bMx8qQtW7RHNVEXBsEk0q
865rCAlrC7uj53BAzd2M0i7P96EWz6+orMEd/faWztqWU+3iNHyX8J9P4ciNW6R9Sc7nr/jlFDxA
g8VVvxhhrp1pHNdOlO/vpDGanaHvx1ozwsJPkRnZ9GLpfPdtoKhnDP1PAc+xS49FR23pSWgJN1ax
NMZhCxOO5HfTWpqYlC6/2tI3MNwB9BNUAKZa+A/jID9fLQNQ9hO3lJ6LtO+XuYqMoZ3pXeJQzYE3
xmgVifLe8XaPFlB1lq0NrxEYq0ch/zQ9H9/IUI5B503WDX7OjuFSBBe6T2Ef8bfoC+vwdKZZBeWG
Rh8WsHIHj9tMXQAU1wyXrazVoibHXmGyhY+sFjjAvT+j8QpMsoevEFzOLSPsjelBrSaODWbDDCUU
v7hxleU0m7gGd2XgNmoXrsZZpd67xvgmkHbmRY0hFwiPr1UyP6dc2ksIBkAdX7EEhZv8RoVIaKX6
4ZL8cEFYIUwKJoYr7NbeFVikIvZiixnfGcmOsZpz9lDioqbwxiKvMjQ2rCROQh0v2OzxJZPkhu0m
IWcYeJA9QmWNn3RA3cerpYmW7GwiJf8V+RWdkFiXAsbH33HDOHK3NkAM/mFrKvLAplOdIuHzi3An
A22gE7uQzPRInDi7ax8dIWUioX+RJn2MexywJjGnxMvLdxb5/gKjyJitiFX92veuLhkE1mV6tTK1
aBWyUnFwgqAvpuH3DG07aoy+TyupBCY5r1PmUQbUKFIFL5JA9rnmKgToNykc9d+LaTlNtMs8cWnY
rYLVPJygmpI1G0BfXf6YuyUxNW/TF88Htu2Et+NKxRtrKGSjuLRDXom+1+8OyeKhFB85uGb4PCQp
DHJ4n5Z5ZRkqayLQIyeOGt7NxSRBCQ+qUulNVREW9wGw4ZLNOODMlTvA9EnLMMngXV2WUbY2bsV/
F7z1pOP5vmGi+lDvMDfo0tzXFjzo0FiuJ1/Z46S1xtOD/zS+rTTgBNc5RwXysfShdM8Q5QCqs42R
zuw22mpycyO36Fx03WkuvBvyiyPJcIbGfl9QpvtNH2XSwrlHyDtIapbnWB7VzAvvLsGWFW50iR3N
aigKrnJn2weZ75VqkE1CIeJ12Ck/ptYu8blqm1L+NBOtGtEqtFtIzAg2GJjiJ+xaMTBxVgcXeRdS
zsSzkDA0i0HSK3UIJCKFFWIT2fphE5UHXOnj2/Pl5uDuX1uywAYCFqu+kAi1Pm79zO/kws+xCSlr
EiFqJWckQeYqJdrVmisDiZP62/GQU/BWdpRnmA77OfetkxKXQWFC7vBdSDhSHgIEQCD7BLO2N1Bu
WFzXRbegmDSPunfo1h7NjJTxHs9LgS4xyacPNxV34qu93L3suJTKhGKTApLOhqpfwXm/ulS8Qmhg
IgFAG++1GzcCAPtnAhgNa3Q8YN06vufNIOoVBQyS2t04KezVo7N1EvJi7Sj1BJPbiEI6hl7TWufc
dojGzZfLFEkfqi4H/S3oBfDnUoIDtQjW+9O/0Sxkq9mSShr2FYErg9gGsL5OILQYCqzQRwh90B/K
NU/A9ENKzgtho00+4tzUAnQc0iSeJw1gqzsoyid264Sg1O+IGeBtPg6FahnZ1Z2EMFo+WM0Y4TyS
mOMaWpzV2Ij20Y2iUGVBm7Y+vlkZ1MsMBnTNujjqJzLmRgjr3ctlTgd/IvppznM1sWsxN3Z/Uj6r
uWq1x46oEmgRE6KxZpcO3x/WKrMKHZ4xdqjyGLM1hX7blxd0bfCCZar5/EicSwluV1Hi2UGsMAwM
Oe6v6A3h7gMmsW10BSYy4pD6D1kJzXQZxfMEpvJeMTkYEObPKGDJdV9ArQqlGl4qnPLXpDNi9Ujp
zoAYzG7/+MymWkHXsYlT3C75Z0UWbYige81h+yAPFyHzwCYDK3/++/FYEhxmAYC8tYQd9mNkx0RF
4IsMuCgy7ep5r98oUbv6UGinF+F+/hLMoHfD2tmIAF25wO7M9OyTfCRU6bmOOBisHTI8s5nqSu3O
2OGjoPHQ0VpBNNmCDpvsmPL3IqApnDXtQ3Pwyf0vUrTt8Gnq7eYqe2kSZdXjAw3/gmeGGVXLClnk
GHJ/4Bb3cZf8ix4YHJ2SGgtSn71W6um76W//Z67lZJRxgKjOYW/hBqpas5a2QXrh/dMs5w+afofn
cmsIq+tldFu1BzleX2ocDR04ENrgvb5ZTUXZKv0WcdGla/5MN2Hg3/OEN0vTNGDXTDkQQT1f1cwk
YkzJp4o76zvTG/Q/Ao3RCaTwN+4LxtG5j6uDPHJYaNfnBEuJnMAyXhNlkjFrpp/LsXc8nc65Jsn/
uL7cTimp4xpEhoav86ZDKxz3F2nsZYPLyX7TRcOD2yx3MkNEpg4YJ6CbEnz5cuYQZsxJSbOuH59b
sKHQjI5OrF6HXvAr4+eTrq+VkWLAain6jVNaiOn5FtjZR6yxADxDGBgWvanES8QikeE73lj4lggJ
fCvzbb4ZeLAjPr7IsqjiYORm6sb83tqakRDcSaIGXSQePrs6qYt0z2JZhbxGhjSOC7gzrg4nYXm4
Udj36OCrQwwifsVHI+gQWPkwv9DJNJk+sT53BTxWGr/B31Oiiplp2iS7qtz1/jEQ+dJyKie6Tb8Y
Gw8kiMyE9lSlxAcFoNZB1b69A4e/mOwgPrqIDKXB4TGDGh+NVrGAeqSOpYoCeq/Ix2mfPeN+Tm6U
44w8UkoN2T9VKin2BK5l/Z3MN9VFduhhDrgkkFmiolc+PlqPRAnHyvjVqVo+WaHKrX4csyIcmVBG
oeRBBza1Sh78h6wkGRuBQPXibMWIRQfzweEMxr52JQ1rGntBvRoQi8JT3NJpoVYy+BgJyAYNHDXl
efkV4H4ybmWELSLiuSiElpxrTnwJ5XN2iiCarpRcfRYZ4L3669MM3NujoLLc2PwYk57SiDW54wgR
C4ikPCV23wbypsVRCTAM8OHi4EFUl8DRe4ZHta965G5LsdiQ55V+8i0USnE79e2XYJCnDf8HNEp/
rXuBOq+Qx4Xh/qJPa66luaX0doUGHzLXaIKCEu6S1g/QjZ9qLsAXbtRWlJMfYAnfGby7UKIoFLEf
wqlqk/lo3rFUaQlVbOiL22r4DI2n9SszUrRT45WiuirC/Lswtm9eHAXm/dwdF3XZ0nRAhlpMtEZc
4h6u67mniVSnAnjacOWBsiaJX8fZB7tCXCRE0Ys/oY9zY24Ax7+WqVgGi1Jl9lV0c9WFR16NXH2h
FhtStH0VAL56/Ae14J/FxSf7L15jj2UJ9KFTv9aUF3sYvYH1Vb9+/gicWB2f4vuHfxHyGR2ZeM7W
iZz+zZ8ZiD791g3t+iFKHOxEdqwKy2FtAAg/eNUeJw/SSvuQwXMeG0pKoN4DnuRpj49Vl8h7jUQI
bTYKI9l68XvVV4konDakXr4omleoXXMuDUp5aA6Y064JznIjujrslgbIxEg/WqwOavljmfa533Pg
NosMSzubhC0nHs96mP20H2Bdn5gOhqnerIKEVXQ9vkzBh3EbdKN9gw2MRmBJOZuGTCDxqNXm7KPb
O+KDfA8Cgf6oy43UftmBuaq9irbE/QTApJf2K1Lyo77hjCgQh2NzVLh0voeZ0UfZW7BJsRODWcNv
va5k8wMdVi+zew4g5W6WQTj90dqVR+bU3vgOcRSIpv4bNzHz9NiXFrU1zIJ7sr7rm5BHevPU067i
LpW+r6NFIjyvSuKSfpqkc+WYpZ8TOWRRkeCbx7jU88U2UkBBos5eCywsUxA979twxGn+1jQ+uTgB
4yI+ocaKfGFKVMSo+iAJYJU5gtbzVFX3f9WwWUL0Jvgqwvb5P/hlg/HSOG9pZaDzYcEvqphOG1xT
ZKTsBL8ieYcfhkrVvixMkNr9vMkG5llmvdlIzwILK9auqYXAZ2aTti/5mBKX8LrQBu0zLn1cDzmp
fuCTKYOmr9N6dUbDHTkdF02kPGNCkh59Rm/zIvn0+VFK66l4p4Vq3ZxoPa39rhXR7thc4ZEiXYh+
7ZrXuxzxPyqyNqAECqGyBamx9USVNBx91h6DNFJ7Kdxr2Xm7D04ZKm3vs74a8MhgSyn4nB4Jm1al
T++2n9WyvtNyLzhSetx/WhnPIhomifgZEe9RACjWGLILZCrD+EssuMDTNXQV5iLVPMvvhN339oev
0C6wWZc4M0YK+DEvPRVDxZx8qvb2pIVffmVYETiiqTdz20GbAdlQH+IDxOF0lB1H4jmno+xuYpH3
wKr1mN2KVIEW7nu8/Qhd5owy6mTuviM3AisTj5Z99sJhhPaRHUPgq6QX+PSJFdFZhgYISevdW6To
zikt7cpCIrsHeJ3d7xLCnZLyX1cxkb4y7q+6xZXOiFmOraBXnsIOYVzH+7lN5Il7ccFMWxmbehcp
x1jj5SU+URP63Tmui5b6NVjUXdJserPQPO6UveBqSc7igzEZ362CcH+222HmbFyVtqYDhXz/iGTk
9WMaQblKJE7Iw61LZjO8HD2P8+3g8D+Vo6kJIgnoBtR6WOTRmzWaY1vHJx0qdBzFDX0oVyeB5fW+
Sjr7eDCQRxTBo6vJ5vCQ3dmLizwMXsMyWJkY8Du7ZaEr3FI4ZdnxABljjDM7cgAxvwrtwgiplyrt
RKmZFmTxVg4O/Guk7t2hkl6mRPK5zs2cu8LEeASORnpdnuIKpVNhMVccX0bt5bnUlIHn4pbrIWyP
t7a9szSb+fB7XgXsi9jJjsOwuN3VBMir7ocL7XARi3a+YJrIEMtCTeA7/V/ns5Zg0rofzhdCKWVt
dVEPtIlCsqF7ekmtiGGtBVMhWSdLQWKYLcpzQz84hSmC0F1e9+/0VN5eM3Qs9/WUJNsf8ywfkECb
S0j62uOGlsctCvQXr/3SYFa3XTld0efBno9uGRypMfBJOX6b2zCi+FlDMZmOw9T4S4IriYrQK9yr
32ttesfWPqTCMZPi3ugIaO1w5kvY7clKW6bpMLp803lg/qvFZt2K28z2X0JkMtpyjdQ+rf/TrgRv
UQDzh0UMoaUd0PUllfd0RbBjdEOZ3CGtFQwNLlj/mUYFMeCAMW4Fee3SWCiVysZIK+sVX++f2I8k
WerpBztx36nRufnrOcsu2uW+4Au+YcMC7dmTrzZRfrFf64ojIV8T5nq6q+8qtGMSGa5eWcrBvULk
9F7aO6Bd21RGgPs6IQO/mhDrespeA2/4psF5mLVUHZqbzrAvaaM0NE6vmt+ar5R0CsVYhk3ZvQ43
USRwH5EJCaUG9hPLBmhtoKN7ulr8ZmHpqDzvwIAW0KOeV1HVKzKluP4KdQWCBYlZTSqWQ4wkBC2u
HRYgBYVQIekvCp/5qY3mwnV4mJ3tcyJDwPlp6rZ5qiLKxDGI+0JbxukhR8SzXy17orApW8WaZqw8
pbU713s/Yca4kKnpIdw2p5TDtOiIOyVAK1b5WreC0nphglq1rcg1ZUvQNrwJdJTHpYEU1wQvi4//
Jp1Uzlpt8BxVGB6+SIO9J2p/XNyJUaj8G33y9ar1A16Agx1EWKaPMYkqAYjXdx/e4WLd6ePEnj/v
T4VNRhW2KEvpJ8h0xqoh/liEwYr2koH6BOK6b+qbE1CUbzkv6HyJEyQN8e1DMyf64xE1g+Vo+yi3
SqdS9iIITW58I7fO0o/ZuC13uUhL2RYm2aC5T8+b7dORQpCfP/AqtvcMApxgYGU+1gpqTwnv90jg
DyYkUwvl+CZqvsMRVc3VULr7/tcXLwXiQp/qXAil78r84Qmuj6jqamdiE6TKNi8kMvmJJcF3XMXI
+X3YZTo0zxm/bT+hf4LhSVepu01ZOW3Cp3aHqZLOBtFvG34065IEhgpjrND/Z98Mh+wAwumZfWiE
eSRIS+Gv/eoht2qLYb25wgn+boX5poPX+JWrkYFktebqaBKkvjhMuwVHFZC47BkW5SkJJ94QkNXC
5vCWrVp7d8i1HomG3PrY/IBvb2NGCKPb3VEGTaTg63qEg6D6VumR9nqSx5RujYZK8YeWMFKJ4YQ3
eCxTg7TRoAdxn9p2xKVFmVbOxt9trnztYWUPIQzx8R1U/ipqx3n5UDwdR3radDZDfS6ICvUbukMl
Lg+1eUfTvoK4fojNcn0nYlTvU76wJVyfVbGBKWhqbBjWszq/IIj4YIaeRpHO/qObTPAbt/FNjWzm
32wOLZ32YXC5qQDQLrIvAqIDNY7dWllyhquGUZjziWSE6THXDUuyy6wWHVbJd4OcKE76FYAeQyZV
34ucz6BEoMNy33fj1baYRZwwOcSBqDmxNv4G2ZF54/0MJRFGT83VeyGrRrm3xpQeInaabRag7LRB
OjpFNgD7gncnZnvjPUg11fMzzbZzT+81MWu4EYzK7wfLBhtmP9eqLL4ioASK+GCo9fi8MDi3KoMr
xx7iAFoL0Z/khOZ7vNvqTmbjgVrmIM2Jkn97B9q7DazTn0hCHT4KdTDTAtYKFpXutzPNKMNu4ZEL
jtd50+nl/ocMPJfElQoDvTs3HFhtiGp4gci3hynB6BgtG8z5UbM0Ihnbf9amg86isJB60MKUH2L+
LN59zskynWVY9PCFx4oy5ldztQqqmZgfBnJBXCaw5WHf6QlwDLVWMRyNjkaCj6snPP5RCABEg6Y0
HcWcB8SBVmreCrT2KtwWQGMGwk2WTgq10WdR6Lfrw2oBfkqV4PmF4IRwtsMOJOIgWeRWKj9jTFJl
4IiNj/JZOWg12arbt4nqsx+D9QMJm6QbYH+Of0DVU0743MkYye71lUAW1Xrwcls8X5sMICz1TtAg
mk7XNL1gZ5bAnw4fF4nWWR6Dz0PH92fl4SJON6PuZ4KO0RnuL1nNjlCGkSlgLLVDOxT5Kc1KJ4rB
ld0RPesKDH35mPhLDdmmk73cJrYeNveViWjCjjK5TeDnHXjBZwDhFFqxFCUSAK/qxhOt+OItDZe6
H/v/fP0pmOwkXhTsU+A9biLSKZ6Ehj5FkN+43bnRfcdZtE0LYzGuWSL0BK3qfuy8bsdgk0zt3F9C
DlrsBSqomqn3BBFRP/3BLXNiAXXTOwiMenYgcSp5WmDjc6r/n1PBZW+/CO/YFOwVm1nIUKrk4FaH
GC100YOadXXPlDA6/vSxrn7AkDDXoXVYlMf8FB0nly1gjC6XlNvIAREhqnomBh+aDfzp/OSOf4OK
9akvArImujQhU90jjDdPR/uEOY2kCZbrstk1MriV+I9RKddHFSNfhW+uRGcpTgvmoTWODGLEthdN
zADIYqtWh39oKj38ZdS8tmfS14A0k6b4kCkP7r2PNlurZ9s8vCnuQgPXeirAHWfEz91AKdGK/sgO
lAyvcqW+QshtHWQ/kbpq7tkDfOIDVBwLTWq0D7TqjdpDIHWtN98F0QYl9oiZF4TFaAgWZgTACmlK
tBe5yyo3OuxrCN2MS8XWrIsqaxW2Y+/wKOUBjpGRlX2mwzcXIgCDeMV+bYKQIkV9YimQI10n9SfN
tfhIcxYvLzkqO7EqMYIKrZzeVLoY3/vLfuHyxfgF0qg6Fz/1blUomcxTZv8u5ml9Kizb08R9oB82
h5qAQysLRQLoZrtUVLwH4N3c/uBZEmIH8cdT9ovxbZjDqdgAtEtlqi0r6Nf0mvF0F2D+E049coVB
ihWFe8hyxIY2qejtkqq3atlPnXzkhLmN5T9IsduP8vM4o4c7lOs+ouzIkk3KiRAm7ZV4mS4J14Xa
Hw5UVZt7oYnZa+adQtvAgjtLlMDMKrkNYlSuRNv1ulZ/SnZU9aTwR4qbNkFKAKxTzjmy7ELVVUxz
7s3gDWukN+jfPbLmskdSb3cP7ugwazNMvy5XuT21uhWahIOqo+gkU2IVsTGheT3O4t3thlCCnecl
keNokNj442eoPe2pNsQDuslKC9DWdGghH3GTOBLT0/kCGiH+b8LKeij63hCcmIfxNk9XxKfrjw3B
4eK5PJqUqSCG1uuAD7LyvnJT6BbDilZBu/aXLBmcsTZm7feQ3q+4jjyANzV0Hvwy8erKpCRZ0E4t
XoOd1EKhBCtCBUSvZgbrvQEUGcOLKhDG6iUEb0CnwHmWAr6crPkAGs0OLzFK537lH1ExapdpTwuu
zmX+Kf+litua9lgIdsbs6ji981YKvOW4EQdxiiKk9UdkxTNjD0+u+4biUb9fK46p3ew8oeo6MuIA
VbuPS5VqGsaArEqwYxYlLEJo1McsvNE5rVwD4Rh0KSU+0Cz7WVXtQOATkW6NBGWLtyhsEaYQhoYs
lo3gjauWslx/s7Gg+pSEpw2OT79aw0g4tBpttIeVeFCU/NxRM1kuiTPN1mkdvL43GHegIukyFRKK
wn/Be2WTjX7O+ZksHaZDcHC7kgzED4qdJyoeMvLQNaqEpwuxuF7k35uI88dwfV+OqDf0S3D/Bkln
/8RAVeddggRE4c4GFGJ7Y1B4KeKAUrvDEwlzuqPXrpjIKKdten6uPbxYRxiWtjMn93qj9v8QVNFp
fCD7ypB0aqtgzGPpKpyZb5O04y9mjDJJatG4VAaUOTzXGebNZ0aIox/W2AwHXItcNt2J7IyaGeT0
JTpSD+0aYr7/TtqDG5LeWdg0U4uIrL293vK0B4QBnip7dubrwmU3RdIvCMUAL3OR15apy934X5tk
VmUQlFzmpha9HqTXhsJbrI4KUOCf0rAvU7J+r9q1WDtGie19oHHLj5AdJapHh+9DUpvp14JdtxVl
eJ7rGkKHH8wLvYLplw9RvHiHaBosktTeAxFBFIMjFqWktZgc6Oe9hCAXQaO9KgdnBWTd4BHTVIeO
uYBhk2qUfay/g0qboBJGKEe3FgwXGU9ThZwJyCQwOhYHEk6pdzyhOibe9MNe9I8dQxui36OeYj1N
dHUH/XoevPlZYHh81/1GOfh8Gk4FFE834cy9FKSkgfP/29sEu1N02RqrhmfCkByiGEeqEbq4AH/b
sxNtAuWRaChhRUGSHRS55Vv6Zc0HtTz67A718HUnX86QeH5UzvuiNR0bDmJrsbGR71GRSE2Ys9N4
Kp2V8qz9xfvLTq+pTOvkBDcwnlAQSwK53g2j67vQVjS3K3x4veD/Kx4O8xwVPy+bm3E5Q9ipf4GB
gKz4G58bbUvveM0gXtnO3yj4bQELuOU2hRSqmWoemuD4EJqg7eXHDRnFsiDsBhj0eQNJEGRKWOFy
COfOA1U+bZJPqP+2nBMTc81iijwxLmmsqeK4kySsjVc8ELLB+I13HuULyAqffZ/8R2tQTg8aKldu
ULDl/tH7Wrzxmhhw3OsKfRHdmO0m8MnBy1ELY+fG57XZNsd42vwpK701cr7HZfJQvp5Kw5VS5dJJ
8sCjc5PQ2/boWVh2chYouo93ILOipEIaa1VbMqhtrM08vccwLKozYWi3pdZKMo///N522jrQB2dO
wATOv4NQrwazxeXEvuPPwO1tNc4HUuLlA7SJvaoSkptZmI5gk3/bPTY8nwfb2D4d39uSq8Y0G/1/
UEz2s2rxmDywSYmDf22EKYgWZgM+eX+mOMg0uQcRxviQx2Dh/KJyi6SOdzkuv5b7EhfMr5PRJR2c
bbdHAyW+FXC+YZ2IPChs10wlJwxg/BZ8pNNWRCBWh8199BbENAxKutW6wRsmJPfuDglADZicmh9+
72Fb05J7KhUGC1Q3t47tkL+7nc6cF4AUmwNzA0Azu4aqVZQrzZ4CMJVkvOOQWJJVACUp+dB2mlVW
zOKv0ZZ9M7NLdicC3lcZOpAeSXpAKqrH2Pu20TdrhJZCEsBOfGUkOom+K2TS3b9Yv3Zikyg0ENEj
4pQQYNScIMkCoZtdfvsGNZlTpyR4aBXA+R3TVFxHcBSWzjSoiKXH+rD8Q/G88MFXb6uUqLEgeZ3Q
iSgLpxvGHpP/Uv1OjuovL/3zDPk7q7WCXsOjnrk1OtPZol6fVcfIvZaOkOcSb3EaoscXWBOIlMNd
qCSySI8TjB7BqY7UKkCXFsgbOtN6IYcd4kR96BleCzkRPBwICXmVA3RXiEghAvH5hgDWC3f51BJI
bgKStw1LxLOfhdX196sWyIL9Mct9IF7oo045nFB6RPpmx1jVIiJsptKPg92p5Vgh+JvbWXn1tJey
Sz1FWVkrh6it14PIL+hOQwdvRhA8BGkfbORUWAcRxHkY4NVjtdqxIj4UGMLhgbe169g8Xpayi9QM
6nyxNcrcUtdU0nXlm+tuN/5nN4S/2nF+YJ3pWM7uP0STtFfe8ON1vlFoOBE3jaOCnnn+HAhRS6F5
JXLlSp/wEngxK7xUsQUBeDJW81R4oPjRScRQT/QFW06CAJMuYfYwMTSKGsDVtcpJ5Km14Gp1KmV3
RyVhO5g3deYD50svWNIA7gxJdBF10BJS/mxNBfjURhnYoAjm+Bt1EAwlABIA5Sh9Jc7SqTx4GUF2
WXdo4F2KJ3JaVz77omPLxlXfTQHm3M7ggjBoAdpYKD4Ce13bFTzW19NEQWhTkyeRpGKGkLZZjfQ7
OAzly3q03vcEACU12fGCYdjPlX/U7xidPKRzxBWRrazRl3K3tz30tkPLiW3Inkpy8z4ATQKK0GN8
vWxcNL2ctvnSKI2nhWHuEwAj9x9K6EV1lCAG9U69lhcIxSBHE0lp/dBAZkQ0rCBtCn2zcs47MdV2
xjetCpxkDG3UarDUtMV7z+QdDm8Og3pVYCdUCd2BXMTsUpCKHIzDCKZUIIojX+2hV3OLhE+bbjiq
jHx6znj960VKROkl9eFQRtaATDItIklzYWuM80VeCRA0Ug/LHwWgxVFDk8f5iAAR50YQuL03DMnJ
9y3336oH5Y20at/oqCXHXqxBKyAiri9D2l0jqKk7HqrkuHPSTTwOy/UMsmEO73dz+lrR4b4Cgpd4
YLB8CEvNc9kip34sfe2/Ki+4feKyLLOAE4M5j+YBh5I1z+EIG0EG2AaHrjoDCTDGpjun7IpBaLEO
jq27TW2jOD8GCIw1I1G/jKW0pmRe645A+G06jMcM58bMMfm6UIEoTABHGpHXhTHzbSwiMNPKpTZz
ArBUtJMs64Gj4nCqKY0u0FSgrbswv8+8qOc+SnRvUFFY9l4j7geKxtD1OSBn+49XPFhaQN0LGOR3
wAm40Olx6tzfCDbpRZ/oo5IvLoSsvyD/95RibLY337OxRZ1o02RqUNivkUY0L2p0rvax5h2eADcz
getbUHVWEIZokX8ns09Oq/qVoNWnGIipHNAseccBr6WAkVrZhxZFrSxvjSGL8J0zAKnzbhXBqCXS
N5jDZNTZMz4Pxc1+RyXuhQHDfigJb9H1c24aknTL0ixYQZWsWqf3cjS4u6y6MwchxzaNfZ0cOThx
f1ho2prCzKxtoQvEtK0o1AV6pLD/jd7w2u92rsEPrPK56VF0F+PSLZKnzDag50w98YqcmmUguKT8
d4Fk8+w1P2vBJOvLylvU9U4OwTMHlF7lu5Ux082h9xOcbBOB6Lxl7OMS1PXyqmVxklnoLrcLjAA8
DKitomsK5zEZHOPMH1MKEENrwrb0YoYPK0QfHKj/e78hH7C/Cf3s4B25twhSMgxJs9yWy3K+DO4h
KoYLlxTKw/rvlY2EI4wk7Z0RnaUjVhBJFI3XirF6/bq+KN6rWDxfgRpMAqQ+J8NpZOehw++7DwG3
Jlo9b7BvHHtcW6sAk9Jmwv1ItnT1UpAhsLxORtTKebQ/FqsZ989nGvZ3VRb1Jxv4tl77hdUnc3LY
tQ8JNiGypaOt3A1GgOx7u/jUfrrtZNh6F43QdxR/m6FLuuoKmBaOSjLuDUB6Ca69yXopoylvgbl2
NYj0bCDWqnK2Ffqn3ne39yl+Tn8uZmLeKDLHotMpULtJ+xBgM0RRKT1sutZYln/vE2pofqEBuibc
98bDlDIrimNaIWkIqg760x5gl83ndIZqmQQf3e1fhUS33Nov4ONj9og+3c23AwpKuNZJPZrZsmf0
yTXxMOITDPKfpm8hp6wekB2HkMcn+al4fHXz4ZB+vulPIvyV9W+hC/CbpuiD05v1ypMtX9XQA/fC
RN+FGpaMvACDfNNFOrXT5VpV6vcQnzXohr88hUoLKzk8XUAnQr9yM8y08VkYG7ZliFTWbl1upyW4
pjQygW9+T3PcNbsYh5uwd0ts1LH5lY2MdxF1dkFF5MgNaB/SsP4wrZVFHcvQKi9QdY/uHt9ArlvQ
pnj80PgtJLWiE/yNsRsgaJo68Ml0mK5acohMH/DtfoMtKZLKYTJgHcajq7WVG1ODHru+UPy+6U4B
Jha/Kk6e4NObje1fS9cJEuVrLcAg27boz2mHYOyHf6qYMEsllneKO4WueJq9DwHBUPAiCCH41eX2
yl4iQ28UVlxWhApBRUYy5evmvnHosmP2j/TXCwi6LPQLoVfHoXm3tD6bOZZoNz2qHht1DX+RZN14
heY6uS2f6fHArrnRRRT5FELBDZ9grM1V8fAYqFjLJLMK5xWs5cDgVMTzMfNMBwQ9MIPHOmjHYeZA
0py1eBtGiMl6RVu9ymATnKb9gOzT2nKsEurVNitJW/jXrXFC+o16+WgrJz4JMGoYm33F3m8f++WP
C+WwtxnBA2xoW7NnsLDV9RNzVr77WOl0G5wkj0dXFdM7poNmlLuSQsZ0Qq2/ah3wSYA5MaP2RGSP
MM0BtLH+B3Ikd9YlC3LMNImc12OlAm9rz8FiCmOJY3wAHGAlE/3KD1QGAJI1+PiSfPh3rP04zUQ5
utjdPqnklThgW4PEZTO93jhhde5YzQIZrYu/yEifWx8Q704uPEMxLcC+zSbAsGBLLaIBs2yNuQjV
eeiprl7exocyt4+IeQYHP2AnxwTa4kJfa/Q5fdaPqMy0Q+BSGW9vvkTjo3J+n/Mmvbq7DILFBLLC
Z+BL4ZdGqyyGE1X3DK7RTPu0SAidOtjqdw0XDHpNycHKpdqDegKkQKb9GMELMkeV1mHe2Oq/XzZE
r5t2oe/wX538yxc+tqnvn2IL55C60t9qrmiDdfiRKerZcfIN1rjqOlJo3drE/+qIeTssCsf6DFRV
0Xhjbgg2/nAxdkYaX4JEq9JfNDP1jcJFD4i3odu904xutGednHtkGA3yLd6+OoDVWGx8aZElybdN
kqarJR3IRgAhZ238JS0sUrCDyX4N6gF4NtZtXu3/lLTw2mj0X1bTm28cdwf0X1cHvSGcWxiHH1YX
sucNGDvVd87FrvrkqrT/g74qpRW/YodKhkuj7FIt88Etsb+eODN60eK1IjkNR1bBGir3WKqubqkE
6c5t1AMAzixMH7OY2IbQ2NgBtHNeg3O3Bw4BGckq8cZjCNair4lQGOeoCp2ISIN6yWLSvG5s5yrM
D/r4AlLGn1G869EKnmDXPv1nJGzLD5XgJVOCnyp24ckgoWe0pDSlLHOoKKepqZRXCurnBJPLcl+o
fSjzZrNAwqcB+R8iojA6qpqIWtbH3OSoI98wdP9A+zsQ4BzhOdSrp2ffMB52Tys7URZ05gIzrInM
4gdY7bhXw7b69PHbEmHwZyAYv8/trBfmEMKcbFicEBcGS3IU/VHvGSQVHejhDdccvs654UyOmO/G
cvSLfHAi672+SqiTusFzdKr95GCJfsEG7jjjuqlM8xoeuvF3GKxbEhSi4ufQnlXMl9G7qt4ozqlN
6da5OS1nwAjPktfURAfStVN+hs/k3CLh8jcMlodODuSfUvNqsMGqHyrdQQyXZcgcDepviow6AXD2
/tuKdl8/WQGz/kUfdrMIguSCRr4Oh/0NuGmRy3PsIaxU2OLJiUCGGnUfJUQzL7TJSmmOj0xykOog
EVxtCsI4RDoukb1m7YCCsYB41u9wDQgkZYNK02ADcF5O8wMr7X0kWhMdsSTffGexemq/M7UwiF/L
J1f9pDhto+OGCw1CzYYJ7TQ7WLZKgdRlxzFdOTff94vTXa1kU/bX7RXbKJ0rvl1O6eRpcn6hkz1o
t+aT0nRUlmeIP/STWdRvQpYYcfL/fkZFMuYjWIqLmf3sB0qQvsUKYDF8ckElONr7M++QqRN0F23p
bXd8reFdOpqt6aEdyP0Nx0De+HK6Vg5mgZpmlDmODD6IEUkMepP8qRW42ytMzBRfgGqklxNRSTWV
daJPIcTjwf/SeIIcBFffVcQyLBkKoKoKOyjZavhLnjHA2y/I059vRrTUzsz7EikMIjDMmK/4jUft
ZRCvBLsgxP+75sTFF3rF3uaaBq3d8YZPVPA85EA79R/C+FVkbx4rTTNzJQmvy/+Bchpxyn5vOHta
MiDcWt9V7M1fWAQxMDvOcs4/yeSXWWRMRz/CESq+5bL2zLjhdEPXbFV6nZ/XDd36Zq++U+fBKSEp
NutVilb24u1E+Ogby2n5NsJmu5R1x0u7DoBdTDvRTewZLwRI3CcY2UGFDQqr5g/6uUJUnrU7KdF5
6KcJV5KuczVeukFVJcscMnwZGMwOpyCNWODvCc2sE5oBRSX3IIU+9a4Da/uT4jhEBUWGUyUf1E1a
QmjpbeX4Y1eQrJ2yi3OLxahcB2av2YYdicFjw/zA8inThn6V0PrAf9E04rmCRsmUOCdsPyJ6xXyY
S9aiAgb1MOjmbGquUyoG8XN8Kib3GRh2hx8tC0rY1WEhwn5fT+GGr/3MjYxxlu73cOyUioM3If4h
VyQiri65tKAUuFKmfOFt7IlEDD3tom545SHEr2l5DLiwFP0PMmaeT3+AtRJ/I9Z4dlutWMV5bmmK
AHPOGuomwHMed8tcpcMZm3B/KB9d9IaRii+c8Yo6cjxbzXm3P/9zJCV/eHtShUJYJ7ySE8r4IlRk
ZpGCUhljYUuoS2IfwGzOempCWLo2OXEOt4piL56iIqrLh3wP8ePtXuhO+LWcJxDPBcNzJd3BQEWY
GK3ySHhUYDUG/g7hXY+0Ls+hf/XWrDORBaXQKfnunwEhCxbrIixIS5/+crp0dKP+5Mh/Qx8oKxXm
e4vP9B425GL0O9aRDq6qlX2xeJeOdqrsSD1JWD/1YHBdHUNF4yOh6lpmvBp3gAhU43ICC6UlnbGd
EQ5jNV3ErMGBlzQfGDrXQEtNbbm9yiIdRNLBVk6ZelR5dRdvNGkbgTgHc58oBBzKh3g6GTF/UeNP
m3RVspajdJTuBKJhHTYTly3Hxu25si/Q94CUS5dFkSRmZc/fynj7g3T7hfTc/l1Kjg2B5kAob4ZM
vwKuIbReR+Azfitt5+so7Bih9PBNV1NO9vRUBdV+mYVqAAYZRrpORHgEC2wWWe/k8IJAnM+8gjnS
GhsEkkZYruflZ2ffz9WxxuEtOEqNz3vTTAy6OsPxOqP4ffBoZ1AkeF8O3HVGsBVytscGe5gthxpz
kxptib9WA6Eq5d+nh/kxbsWtTTIDwHid0XNIR44euilVQg0Y3bFTKNO45LVIuKYJCxrjOwIJuUWW
S07D/Jy0QnZx+6b8bsjZbUs06WvUIDWIZSadaLBWWIS7IEKJngtHcVC8W5+LLcmXlxOweAHBUdMU
PPm5nfSc1puYFsbk4RfcVjRHs4TUPMyjEm0WrNsCYVfoAQ/VT3syPgXD0CNe3AWGsCYKQP2Dfvir
/Nn+zWVEub1jNwoVMf6QtyXUJxEnBbupDox0dN+0Fqx2NuAK441MC1P7LKB8KIFLBY8ifbq1KSeN
N77KwkKlLr/xSn2dF2UEDAtBNG30gFFc+WCyR+9JVwCE0Te0uqV9h4BmNbaxitwUX748tDpZVNem
zXeh06ZGUuskrHt9hkizThCaA/e9jQGRjIEDPklF2TFwWlDN0gzV7JkNudI/u8HXVnYZz7ie6cs+
h6/UgGuT/D/NWG66x3vrZla/ZWKnk6KNElpQbnuF1c/8tcpuGR7qoJ2aa5RBG6Ag791AecuByyUR
gqcKJB/z4rZjwu1PlB2gqHBVNOPImelgyaDsV5RHVq0hoe/kgevp2RAjSDmnlWxW7UKRbtYEGszn
3/puhnNkYcG92UWfB5JLFOYcWzgNybZ3X6DX4yD3PimK6ZqaF5qebyZitbv74IN3ZAh8ql5tHk9b
7y0ov/Pj/YGi85PDarQ/oq3ztupHETCsXcb0beFALn86hrj0tjww9GnndwpEFiZfR9Mxsft9mNx4
T9Vr/pqoNW3U5pPOQ99cMZXIXxjouQmXcV8QxauS2exz6NBqXjwSzc//vEOXeeROyNOC1ezqnmLW
O/6pzQuF3WSWU3y6/uKWK8oSQNPbo++6xDnwmoq8IGwnP0bldZXhg2LSVjXO9vhXm6A5vkHe2ZPG
evkNDaUHXKR8gBqX9pgs/vPj7JAmoOrXFJuwO6Jf683GVIcrcnyuaOzRHSp599jqJcG2CkZAlowt
Hzqh73ez9skhBZ3GNAwHXtDVO9/6KGVXXmVzR4ZYyVGDMp4BwiC7ncZpvNLNq7RWoBg5PCo28bD1
jHZBPXjMlz/kJJJnyTqO8Gxc/g34nx8eVwY86zvRrFhtmoGe3FFXe4Lg3Ix8rx4x5xoLzJgunL+q
8WIP31mV2I5Mjb93mgV/s2fIU27qnzBuBCwk7BPFpYycptBzdXWsWy38vurX5JmMQ/899y+UjnuD
tHFWR4nRDb9cH6XBKdwGHFzr75DbFdXhf9NPz5gZCMx80F02o0Jky9GitMeUj2E6icYxVi7aCYdv
8nCRobjt8ZCYraqyjigE6bBeUC6uZekO8sZXFwUfirXZtEXVSrqAtav3s2WDUZ+/KGHRnLIkQry2
ECc0hwAw4IabU1VD81OuqqHrYhAkz6NHe1Vqv0P7TpSbIOx/wexr5fsPB/DH7mKydimYP8lHOOyT
XneMJwTDr9ZSe7PGPDIOObsRuf619HlbSOtkMCvs2b5GlsmH2l/JPBhfBFha74a1AWk20Kc80rrh
EggdmGAnYVsqA4X57p0WFP2h6pe2Q9iWSY0DBFNzUWjpPqt+JQJiScOh0ko9MitGWPhhJf4a3a2h
fx3kZF2e668BVMDV968b0ArRsQgP70zWLR4GBfkPSU3+yNWtXL4z1+3ueaoQDFuHyzBXKBM2lUYV
wV346QyzOaYeasBtMcDpkGIBgYqZq38/w6HftBEpSjKkGocmxvmiWHvvzFzAjq9K4/lLY43f3AJj
2OBoWgfaWdl4wTexars7elQk6ahX1G91tVmP1QMJQty88kMj55Ayq+8sXY8YYmS46+7J9zXwsNBV
hH6Jcgh30DcnWIFpEnlsEA02yCdmvaDPpRS7bLncS3qZWa43yKdqqPEUN21owNg8jOlSx0kaoR8k
HV2JkA9v+tjMF/XINAiQyfEp7jMm2mLpWceJP0vSIo2qSKO8N+RLqHR9g7lyjG4rdLIyCD1uZAJy
Zhkox2DbFAN8oWjNoHnurgift4W460OHLQ82dLXw9lV6ILcqyEScEAQSOLlOuesbdxnHxoGzz8JR
bXz9jhapHu5Y2OEsVwRHBmd2cR50R/ACGv5wAuZNej81gvJnmNrQQHeKZGpzqE215Gi7tdu65l8C
0oA1ldwE68H7O/H89+g+tMsGvy+SZI0J6RWNt+sGZTEQhKmkSny16/9hBAZg89jDb6oBHvMg5y+h
5wBWz6jegsQxH1wPZIONuC1m5kBf+VbhL3iPO5KjmGPeEXbSuSpjJJwQErtlENamGX3CQZ+ceLvg
EddbDYyWREcxh2o4SyDZHEhrNkh2is7igWFo0I9SXJFVIzAnoM4iydlwmZR2ggiltCx2mVPQBgyf
t6rVN8/SXf9zz530o5iKGQpazUBXVVyjVZBtYpK4eu8y/yfNUOAFXVMMzWsRpfZBcXBH57SSk/E5
71R8bVKG4eprO4USq/MZt27EE+iR3g7jLnNzitWc7ypHv2D276rhYywZhEA3KflBCXFYzxiXBalC
HVH1aBNXRQR2zRP3Q4OSxdMWQwyXdyI8UmLFPPJQBMigF2LwNHNXS1g+CvSR2ZfSW6he/IVOy4mk
oxHnJs1jTA2Srq/vosg7eiU9+5ZdgVkjvs6IUa0DYm5G/GPr0FcBYl3khgX/nJxl/x8gVPQAa9qd
uihBsdssgb2BIVrXCQGocaFjvNUr0wUYwjG4mREv2AH6ELToUAOhsQoUjkLW9qLReSTjpRqaculM
VVj4TTV58LVKEwaQH67AXWlAQHtd3pcsfQaOMSlWipwMwV2QvKN9CmvriVasst1VJDGCFxRe94nt
N6HpbRhOgI7evIdbqXftRx3qENaFF6pR/rVcqC0xOsbK8K7nMgvVdwit9mBevRb7qVmepzR1tPji
eOGmWRu5978f78IUt052yZ9crlt7tZv6WrFTFY43Va8pZd/eTQeOGwnr6pTd2VoGCRiN4JJl2ssC
yzdK2OzQJF79YdtnBP9rQUhStwfewp+kV/Fq9rJxL4OvfRUaiVfblCgV9dC5zj+VMvecGonL37l0
uUodiiyib+wRg6NuPbK3fdZnfmosK+S6UB7qH1W4US1zd+yuzNkwSLSfjL/TZ0gQsbIxAoylNR/R
kjhXbHhvPWJKihNgsp+WOdiyQiCI9ctcQ1bM/83gwOt4PVwaFxCixUuMFTj8Rt8ZDqzbe8cf7FbM
GXRz6yY3ggIiMW6s5yiCJyK+Klv/rN84jhT0kOmCv5v8RmuBbpdTVd0CwU2JvX2h+99jw3QOWelG
RONKE9vZyhcKm9XEPAyfVvKX9PhKZbi3cEs0JZoC67HMms14HuzHLk4NyLaaThVFbQhe1ladrrAs
o6VjZkvCo6luVttpCN9/XVmbKcpriWCNFEHpdJhXNqjHiNx8N8dk4JqSSWAyq3toe3hUBT04Fq8u
6sAKmBrZptp4SUM1eArUnFEThllJpvxkTdC/e955f2HAKgOFmm8j70CPp3mcTnLS/9FTcz5cYr06
hEpugEkDTmL9avzU1t5WcboB3hhE/JHRiyw9fzZATRXBY4MHlHQvhz9dCHzvkD+ZqoaLRtEAIgWD
XmIqaMTwgwZbqWno2EdE3axmxFczukOLWY+mn25CyJyrCwZDhGT6qMVYjUkfNABTl0R6Go4AeZxa
XgfY4i1A1/JRGfUSV1pNUXAZY7qg60v1at2BxEiIiqHd2UK0VXD015T7NEDk0qM8LuMCbjgsbY70
NatTkS/iQI6bMOhruhmmmiN3WauGzp41/I7OQes9Q6nXr20qzr3OdhtKWIKGdKiaV1kwDOqroevm
QeSLrjV10ukPub9YSAlM8Wyq6hiWk1u3VwLYx+ovl5bTcN/DAiZ+RNIwl9ERLaL0w0WYvlSOTHsV
RaL4D7c1xqdevy3/sh9Ja97+htxYGSUKN1c6eU53I9mPxP2y7NBLNR4861QjIFeZ255OowoK8qoM
5/0rL4K4tZSyZq8ymKNUixCWhrd+TIOXpGJCGsuXFFM1zxyy9dBvXq8t7u2y2l3JFijHM0BroLLC
wvsdE1Q41GOvTkkAvFl4jGk87s/VT0Sscgaaigq48IDgyq4+gENFsL2igA3RBwl9yO7FSzmHngpH
0z1f1Pwi3rkbBjGsro4AEn8JZRwOzIJ5WJihcYGP/3aLIUAksHfJp5OI2cAHvjReUzIElkbU457Y
gUDisQp8rNF/c6V4/e7qLmneAsa9zRXEQfy+ECtTu0uWbzx8Qv96b4pJra8Ac4t4dMFh3EFh5i6P
1kOmFrTHvwjBMWG0tp/Aj55MPW29K0yLeBuYFkWJW+iUABZ9b71ZSDnXg2LnLngvSdR/4mtSh/R7
ZOyA0BZUJzbIdgjEjl+BffdTnHqtG8a6ijpmcgdN0zo0Peko4hRLW687az3HtLwK63DEVYHvF6a3
E37/uTkTZlqmIx6eUSg+UyyGDXYuDvUs47cUKeqPy+HAEtFILz2O/cTJYxeEK6UqKz14g6Cmkwux
ClfjoQDo2bRcWjq9XvGGhGR1FQLwKjdDiMsv6cNUuttd2x81NYXoSNzot/CUwkaYQJyN1Gvte6Ae
ljGDDU7pOHlzt3ymD/HQFvYScX8Q7+JsZQkypndz9xsiDIfF8o0atBv7vGDxt539vztpVXke3j1J
tay4lqSPhTJ2yYrXPLG+1f0TsmCMrc+LFvn3Cjn6oLw1uN/oYedgMmrn59CbjTOd1z9/qobBInZQ
bS9DvwchAgpejh4Dng7Re+wc5pYsf6vfexIYHb8UU9W1EBmuoAIdzmh2vjrR3uATIXyPyq2vCtWc
HB65sy2r1THU8UhruWZrwO0Or/1B73JYBc7qOSWYLeWhcCX8d7c5pYl6VyzFH9VVqPtMitt4hUcm
eecEXUROFsf7a3VjPA5JSjCXXZM+Gj5xsi4/bF0M7ZY2CVONf4+T612GWOFRfaUdhEdQX46DmVqF
LI4Io/ie6nB4TMQnLCi4mmfbHv9IH0B1pKiQg19L9P8spcWfSaJE00BTsvDmZLJ533NP0s56cPZq
hQ0ymX3dOlWKasZSNx+wDJgf/rG7fvd/Z8PCzwuM7r5yNeDwG2uprA9peLdfB+ntg457BNLFcGBw
+fHCUSy00BxQ24FCFvW5DN/4MlJHsAAjW+6x2etySSgJlbSbObCGAE3+hQHdYdOyVBrlIsiEgV9J
zPva4/agg63nTwyfWHnxC3kCkY15X2/Pgv+3bzwwcd1E81tj9GQRZU1TrMEACX/VH999xuqZo1I7
BOeVBVLo1ByO8JwdUAFsaNGtrEQKQ36hvO7ez2vU+WXbjuXoxEg54fdRVtSJbjHdvnwXlnJjp6QM
hZetrCyDjXInCXZNagVhX3zx9eteyoJx2GE9ZaDJsJ/IOj8mT9Krn0qbSVe9BALGmsv4ci2hfgBs
Javt4QdGXhAGyleZ9IkfSXCWyP6Hx1cjqt6Tl0suwUIaLN+6gcSAnnTN/eknOXKFdwjmhrPtzdzx
sfvYRa+P2Nzj5FXvmVRfqhj8ESuuIXi87BPei3lDZWmm9rWmbIC4Y1HdmLwHjFj7kT1o4YyKB6wq
1DRgwSCrHRqPFTjZfCt36cC87kBhklHc1LVgmuYc34B6M0B7VvtZatBJNznU1+FLUjrwmPTeetBe
3sigS69aWUDH19bEc0JmoyfOIgofxakL57AQHd6lWp1un2F4/pTA/pHlCXtsEawM7DjGsYwucqK6
UMo3OBTURjVlmJGqCBjeFGoDPVEqLjQ+VBymNolHcx2g2OMW2JF9k1wrZNsh9SJrndgTz5hI2okx
QTHBgmxadvqAp78TGTLODYlQebto8Plxwj2aebZWHnoSMIAgcPFgR3PmRbgT9hhkykA78M1SMXMF
aMcW2IQ5yNJxzBmikdncQGe1haMVUaqRyBD6O8Dv+BJI7lO4c7I+iDllHrrpkK3TieK+fzfnGVjt
yHnNMvafmgIGm84AHqByPeOLbYgadW1sE0z4srQSkG1X50EG4L8gaMV+OBmdi9VyOrhIY30mq8gj
XB/80vhub3MRa4V43x8yjMB40t0Rwuql+uw4GaJpKww47uQ5vtImPDyq/nEBjIGYYv8DXT5exEON
God+f2fSND0WpFGYQIQfgW77IGSFCPcv0EmYOOo6k5BWhGsYPE3Q/Gr+vNzfFAL7BCBvCRDYMpCG
zL1mYy4df/Z1pietOpgFDlqaNGiFwthnALyBZt09AWOKLAF8/6erKiFF50x6QwLngqxBgh5D7KAE
vQsRLIVsZUm+Zcd+5kxH4uvyVht9rdPcUMtLhmLfwBJmf9vpngZI+XBrK1mC9zrWLKuGnAWOt5g8
JA1mGjYAywJE1bkSgumzna50oBuoYn4lmCt9Cfipb3GGpSYa55R6KBjmaOJBHPbW8EMNl1dzLET/
em8KCOCv2S89x8kPEt7XsLUoFxcg5LTNRNDzcwvwBwMn0wlJ05fQOOLJdsDb9nVB3+iuF1jzhtJe
9Ma6JV5t1IDlA6cmv3ryA/JFvuX1FsUp6XjHJiW9GvVAV3LwrwAghV+q/MPv2RjXzNRIPVxI3HK7
HY+B3O1VFG0Qqo5djyJ2zIYDEd1Nc4Ldro1XwcgIVGKs1LHY5BXQJnizI5STWwW/cfWWMIZdUtSn
pmEmQWrlzbGwW8PYO0QoD6rbie0ELCSfn0u0OyhIp4/mdW2Tg5muA3W5fICWoBZTF8cAibcZrJdr
weuy4mlrmQLn0EK1XWvtm4aAddyhXhak+R7DIn1iCEcgy9zMYhfr0H/BJ+bbubEpzJGhfbngZD8Z
rkhyqntADrdQCtdHLS8agPvchUs/BELHR6+1c0I6U1n4UkvDLwUtvDDBZwaenHBlyqE4izVJj+XO
mjcdLe6zCLRmJGD3+iJCbG+X6bABaSkrfZKZYRgs/WnJcjVPtCxdSw5/J1lRzcqrJz0IM1002YHT
WBGz7e6zLl+cMnuDKeAL8iJ0xn1ALLt8Lmsfu+rEGvkKCmpVhTcR0S7HeSRliHUu/Pd/Xx0vki8j
xanpt04lZsrsjf8ft+y5yFuXMjoY97gHsaoA1U4Pn4BtKmR8YnVGy02wSlpImJxmbgElRKqkk2aN
YfF/bBIgT77rvRqDbA+5Zvop29b+ILTV5cDSRyZ7oZAyM7t0EghizCwQJLv+t6Lc+BeqTXXEoiVZ
wVeDf7z+MG1PY/vHJKZRRrSpyUG95jmCTB5+0lWdkizmpr/vPeW7hnzpA1WFNk4bLmtNOlD7nkPW
hLZUEziaxh1HoVyd8St+I52J0679GAgRFPXyqIbxXfctpb7oB9qWACr7y44QdMX1Dc7P1ok0VocC
SjEh32EhRg9KJ35l16/Ad5j2gNjboEE09HbCVsmsC0lxmotJ3HTApdCP8VB2KS123O/bWIu6aC7h
XQl3Am9EBWkPqTUiPkXtwIdYNhfMmg0KD3mERy3G/8GL/aVGZcdui8/O8ot2p2swW7O4HsBb1gL8
yiXAY8jXV3feymklWSecNXvMb4JPs2cYsSWqnxwhmAv0xbxTLto+B9ZGNlb7beT64o/NF/krGurL
0sQw3bhagf2mufmio+DO8GRe3r9hWLFVEECW2MRDSUw1deEWs8gT7O2Tqtr9Z27fZoSKn7KsE1M9
J4W34F2vwTd2Pg+7Kbq8ABd+MdtVgZhW5ey4DNfZMRP8itqCfW1QPjbAog6pHnS5/lopyYzVOmWd
ldkGUZ2VN9xD04NgMCwbcJ6NKaksKR5iIwx9Fvo5kUi/WklnADMlXJGDOgnDeHEQtWidxYVvf8Ff
V0asLJdCnZIL6Eo1qJgcUFyr/beT96MFq8VqqIrE+ab09EFVc5Jp6YXK2P3+b9LDP0m6OLC9SbjY
1iAIL4ZDir8PPxO2rHMIUBhVOfJslA2y8zvzCVo2cP0kZTHeudWiY5RCPgiKOPgwQ9ABcxKL2HG9
DJIzx/Gm0QVEBrqLD5P8UtU0jkwtsgHhq6zUZ/YXw6ibnW+MqphbTXbotNVqh5lowGP6zucjeX/d
YMXetmQCMxk+zOMx2e+DpGBZqDbg0caUc07/K0r3UbabmijdGVaUF37vZEPZ2mkk4kbV9x9csK1b
odYzgZt7WNXlxjy4HXhuFcX5NWWIDYxz7YpO2wCV2rxtwVou7zNTVH3HxPozetAvdausLKibkwpk
I2+KFdCtEhKFBGe95XCoNsQ5UnizEuOCAn42TKAc116XuNJO845u6CLA1ExhzLlaI4U3fjaxcHYF
mviCmue7ES9orF75T4DHuFjQPsGsPBwq07k37PUV396RfKSHeXsMad12pkoMfORRXOHUDKKQcgmI
Bo7ToVF0N8DowDeI8oNG1ZfI9RM42Y1I+KxjRWs/o4M7TkVf/coKuLaqkZ8vkAz094wyqenTSb7d
l2VAMaChRoQlRX+KZPah1CVXz3b0FA2xmeTL+zPgklAW4HP15scNCxKDoHpfK/d8SJo8MeEtICtn
E4kuqgaRe3IoLAhcTeR35pei3wuPyNlz3gCelSVuNARtZI9QozwsujtPv/EvY8ySm0Yq0waTm83M
HhZn0n4Q7QTTIu4mwuIE4LQk62OMJpRWfkOp7bm2o7hcXSn0staC9Cr/bOxRZvFhoNiR+B/53TQ+
UEdA7Q9gYp6z3q1RUZnKf/gQT0S2CtGCygTpW1O/HIiJBnr8TSCQwLrbU0uxRB9q4A78S3vYRdIQ
GfvJtyNGVV9G1K8/nHB2ZbtMyJvOfno87SFGN31oGBvdUdmKHqjcXiJaC17SGE35JTbs4FQo5oaI
9j7Q9WoJ3HGg/eXvAWOEwkIrjpfXZol4DYVMECuDL1+SvmtI0wEKnCEQHTENlEbNHBiq+Pl2bPi+
jjm8Ubp4uvFOEVw+EjXcmPilJCUpB5rccDWKXaUik6Q5JcUQ/n56+5pwMvZBehL6kl5XUx3yorvB
E0mUxbrGwFwFV6uS0efUPrZqDuFW8SizxcEbX4e3kx1K5FYg9blZ+wV0upKWL2Tb48266w+nQ5Vz
rUEqWUEHDE7+iUMzu9TG2TeOyZ/Yv7iGP8j+APBkoi2VGD4ZghO2Leh6G3By1P8ResEw/Zx/6y+g
Sl6eGLRzOhnxRWILot9JwWxo5VSc9CFcQ89p2XWnuL1Dqv84I53UeTaeECSrANauCUb7h19o0GWx
5SWK/J19Ke/WnmEhqZUjveyPSEOUrKEulXCMfkJhSTJfB/IWiQjEZHrn7JhwvW0OW73DUj0a4AuH
0BcMboZZvSQ9JxOV/ssZp4WzT90VNQaOpvJ2kFuV7U2/2kEmPNoRn+XabrJlvptCt2pqy3gN4N2b
LMl1+RwbJSYlc/THzGefdGmOTXS39g6U+/KLgBT6OsLksgxJnr0pZp/32Gd6S33rRdy0Q2Ni3F49
fYgyK8HFUuES/z9w4FDeHet09PDSsd3W47OaLE0uk8q63slrShAMKoV7wgj5UnF5MgK0pRvUsIqL
HwPumTa9ZSQSoH+lmCwrfD4g2qxN+AhULv9423FceyVWzKBd58uRO5lEBAF02OvS7em+EL96GDs/
VMP5DfxxFI8Xgalq0ibpihq5kqEfTq/0SJkJWxJfOpaz8QZdHbOjRcUSbkvy/KzE7l2cqoikOuqW
5WwTQCQDLLkQJEvJ+LvTtRvLPCTPEDrRVT4tHvZbOYcZWLND/bqLxdL6XkwvGJjRWsAOr/etPl5X
Vd5uLSGa0p0shErlNlpeDYpnQK0BVsjTb4uUebV3hiltYE4D9jCq8yZ9Z8gEJI4OXRrCyrr+BRoO
zZKde3Z1/Dx9XItxloBCQvzBj9jhUZRPQ8t7AjPCh3AtT0kC5I1OBjV/GdC/JYybxF8nLf7rkL5Q
3jKQ+YfnGc7RB1YFI7klqzIiNYFAh+vHfrLDIATG+Rd3U6L21YgR7IK74NdpCMghF2xzPHEta8Z4
yXt+hgjJaclyy2ODt+wxAz8+fTC2Z0HoRys4mzGpIPSC3FerS6p9T6VNYajI9keH0K4YW1mBksdx
AdzDS3XLUnaNGYa9WHHOqDQrasUk4aRd3gtvXA4bWXE7E32v6WGlnMyBStbuc5/qK36b1z6cNsjM
xX64QkfwoLNNkBljCsawdI+bzGzQDabgD5fxys90Rsc03E5J4epoPotjfy+bpkVaAyLN/wuhpdxg
KOsZrlWw4/tUMhMVwhwdS4nXw3+hb933pJ5lBiBo8OXQEtIEa7c3BHX73yVp8WDFSkMrLgJ1SX13
xdQaE3sckbgd6qkF5HpcDFbwtfg/jXBwi+QCI0OBlLkRkIuBugRnql59sqFlPEABHQnq+yedqvcF
tE7P6K0PGMdM9/M+5T6I12v3cDDIcU+nDCm8Eyks2jkdlWfch9of6JLzbWbwvun5uAxFmtnmDuMk
HHJ1qzvfKMjvXxMpzOArIKPG9M795LpWKrZZ+u/+iAcL/e0pThDs3gdUHeQxypDXuq8CLQeKm3Pk
BlcQU9CCBxkM3iQ3zlvB5RnhS3nMOlfFx4lP0vg0ZR9jRXFb1dJnOdFyPpWRcPubhfEjYyX+ec8d
DKYLTiDEuc99ji6/xIdZXsN0kFZyniqHOj2+j1CccNoSA/TNMRDls8GvykHaCLP4aWse4rQKc0oX
zA45NUkpU9yxHsuYZzEyQjINjQPXApNhFPwS/BScIgHau1YTtUJc1v2CUsBk5qlpid/wMpZqOyMW
+hpxG8ZQwajZ8Wqoto/gXh8vwm2bG4BJRDKE7U9LiYreV/h9XVis2BKSQrxzyyvQl87i9gyeZt0n
98DYu93Koi7lXf9x+OoGfnYZy/qbnIatRO/GuxD7DgA6ZSP/n8AFLI10IwR4vbnWgqBGyIr6iXgU
gHK1eanCnHQIJhdtsRhahAiEcApqEpb+a4sMszzMW//Sdx8hopw2DlifwBRFdtUtOlY/siXRncVo
BcqZly+IH0otkFzsepkW3RV3jUc5UGAkWT5mjlatzPkUtj6DRP05hJmHjsPDEV9QEgCS8HCUVN5f
QFFmKSVjquQ2XnYKg28yV5aKD5Y7jBMzVYRURrkfmzeBpbxrUz177Nco1YZf8BPyJpWVzazoqCq3
gqpHne7kyScDBcPBd5kFwqiNxJLJH50CmZkGA55QrMo55KOT8FSw5s3e3L6dfQLbQ0RWs1gP/NwU
YUiN63ga3EFIR+WQS3ALR7kPERuK8uz9wPyLxUtJjEAgF5NirTBFEf6KBxQfANAgaXMpjVDvU+eJ
uSVS9yPxClKPNVB4PLppugd0wIfJc3uOenrUvO/RLsh2WE4AGrJ9xc0HhpRalU80pgiVzc7rGhtq
QI+ZbthIzFcRiJ09jiTMVoDQv9DfDJDkwEL9DhMFJliSyCFse3vKpWBvUVmDA4RnhjDx283XpkQ5
YhEKMmMD4CgKO8X5zc3MmHDvpBKIWSWYzFwcQrJ9HnJhE9MWjNgd64Rvy1U1J9KHCnCSvuXTqIts
nKkEGl/oxsPAIqjwAlGPepNlpEIN3woZEv9X/vkOUgH11h6tiNZTpXcZ2EXfvEJGk6XmtW7K8RG+
BEqg9r0p5hx7c1uCMuFHzz/Oe9t7QFyBUgqPF8nBXBkNb5SfG16zivUCX9DeSotTt9dgOFLsPASr
Ov8o5LFMdOFiQvg0SXvINDCXdKm6k6U0TFnOU1h+IWuso1krrRC8inRg76TGRC2RLW+a5tIxRioB
pC863t/9BA98SAQV60IB5YNSV5tgHVzGUS5O0Qk39hOam7MfrviIyT1ovePoXf+7rbVKebPE3MlW
vz5SlhFj02KNO/zwsy9vCX6T5PPSd/fiwAN5gu9bNbFcDrTmEGdiy76viwlw7mLrGR9XDdhoA0Dy
rBQ5xAW3l6RxIEEyyCFQjgQ9O3sr5mCXxjcB7cvZuqwpDEX1HYi1o4lORX1joZrfQVmb8yacpqpo
Z2StYe9Ucmo8rYPygMOX28hKWaTmC+OVvwWa/rHxMWoeq3Sxb0fYdPdnuwo2VrzvAWackMdUzVbp
fjWI4xVBhg20Mu/zckG9KOW1/rN0PjydU8Ie0rrUUo50+1CW8lavPPEDh9WgUOgamVAJJEBGutLK
hZYeMKuFtLT92NBFV/AgDiwiXz0itr9L2PKLDLjv6m9uz6QkY929p9mjMNLLLMXdy9zRHvPIgQmb
UtOIm+HjUB4fAaM3+0Prf9FgbpLJU+/3gCs27JXMZfgaZe81IN3PONJqGvX7zF2igpagNKsOvqXL
mL2q7HQT57DzA8PA9l+o/xfA6N0yMKw7rloeNu6nVwNEgdeZbQ/7meY9xIwPkElRNh0NIy6COwPj
e/o9pHfNyT79nICl2XJcFq66ITb3y5UKzJtOCO2aN7w6H2r76xE1aJiaQI+qriJMLxxrKA1t+R8Y
ItOPtWTvwJ2GM5ECmsSdfTEx0MtYioyr/crdU6X3LF9+Dk73T4fP3Fa0SgzmMNwjzIGTzAwRDqGP
YNMbetmjYXXNNeVC5kW0pF4IitIMrlkyDJoEcgyaXTWsqaJ06PKyln69M6MakuOShaODOE/qipoG
UJn7Uy4JYf/mOatW8o1d9qoLXMUAKUXdcV9fEKG5rJnxg9vWh+kN/g+EUovLmkZ8zC5x2DWNNiSm
Zy1hpr+pjcRpSSDiyLBtcxzT+1GcKNq/qyPCuMPOxVwr0PViRG59x5KkwgEa2aU3wRU1xWAGytvZ
pVjexO1EdiHibWlsYjKzWdB1bpHDKK3JWIWXhBie1NE3ynhBEwnGFnzXEXZfH7jyUF+iu1x6qp6F
vhuHOvlzsnATjl7m6OkNW3AuA4jpUTOcPgXVUVUp5BeDDLzz/4wBNXlB/vaTMViySfSdXzbMKxGD
ni+D4aSwSokiFMyk6xqz9nJ5aYImuMyAryWuojZ3941mPMPDgdh+1OhM93hJAhQlmlOptvUgtrHd
WA3d3KqwXVFw2EgUSyceDQtaQvvH4yaaHNwkEjjbnqrjQL0MClx1bvPtAPET2PktthHjNfGmmKvF
qMouF24QmzC0JwpJ5DcCdLGjBHXZAzDxyJZmSnKy+ZrAxve4nHmNBl8Xb0/zgDmXkSaFNzWhjNbd
m4DEAJteVw0jKjXaBd2qETZo7zvMHAKSpYVttExr90MSXFZgj+eTeCZZagJTXLXO+RhSiePuoLAN
n4VAMUNBN6hpKBjn/cxI4tyswcuk0JIev64vrEE347Hu5/xn4ubRIZifxYFCE98PbVRxHFhHwZ8I
O8ZbduD+3cHik/o0xLDEszsJ6c9fZNLcBZ3e2P5+9st2nKzaIz5QuQPRo5wMlbM9m+2iY13XkNOi
pSYpvlJ0aqe0hjFwHT5HjPBKurpk+/fw00ExOwDFv5UbSxhTcxD/WhJCZ99UQfmISBZ2A+wwem7S
OeTtLvdzUOUXZ2Qo5AjhsNs7wA3PQLeSntJ0NL24mRHdmM4mRvilvunBQJfIDPeUrKRx9pRiEzyJ
4YvGFTHFSzMV2EDpzChAzWygs+ZfuV/YmBckg/64/gG+g+TyXPOx5/wDv2tehplb34gC4UR2KHkF
4YJ69jfYOXUSagQHia6e7OzxEd7GdqmFWQWx6run08FO+4DQ+PZMsxSNcNIL0mGebP0I9PjS6JHu
lTcD3bk21YP84O3hZKER3ZqrAeQ8TCHrgA8rlBG73jy31xwhZvYyrc9FhDp6gIYj0xjOPlT5Ejab
mMvOjtmEO/7rUeINBH81gMK1vuOSmoktjs1WDGyDUkWyMsVuIi5DtWmHG1HzgI04/ByM7Qz65ryt
Wdww4Y4FSxBhBwi74Eh9z5ZHPJ2zu/ElIdKeH0cnn28ERrdjYo4ljsnT03dLPVE4NhvM8p1DYrJK
BJ0u7gpiGHDaB1BZzGpm+lRctxnqE0bxqIdYAwl2pTSpuNNiGBzMxAQONylvRcpFu8sS0LZR9BgJ
yWEMcVS6MXDMdKPf4LFC7FA0+P5IqPqVWq52MYa0ypDCwtie+rc+hPz9HlAqVULsfNOVLnVunPzu
Id1J68bL/yl9EPfxZjRmLAs4/8yDtUByCLiiqPAWjMsLcsFToKn5bk62eY54uJdAsv5hZE437J7C
QrUnWrNzqCaIz+nL7tYKBRkibKn9JjydTauajU6/NRC2PnKoNF/VBjjck1dsvLyrMQRUVl3Utg2v
xmPmaEs7q4FWEXyioNJ7VS//3TGdYzLUmgpthJSkJDRj9hZK5u3Fo2KSANhDdeJwTgwG1XbgD2mC
dBizSp4y1qHYdLANrOI9HgefyFNV5AkW9aNrTisSKoej3CatZEIUhdwJAZ+t8/T8odeGpyNX0RS6
TMFcyPk/MtqAV987leYkfuaearI0v8XKBrJf54nCIbD1XAq6x1nXjD65DCDszi9+8wWoaP8enEs6
ZlU2VeDju46a9VQaU7ZfhY6ftRjdaDduUErXAEBiWbenFI2WaiQXmXyyWjagHwsqLI9tPiL3g5jU
AmXHBFtOd+rZPIOn0WsYGbpLTBgRdbTAN83MC60APml9DXGTAAjDSwxAOsQzYneQOZPNlqYCWgHy
EoASzX/486dm/bYOyhpXazAVndTC08+j3DK2jzPmTcTyFXcPmagwGwe6BJaQ9vBQKXGwyPXO9VUY
EieiD39TZSINBxupQ4gK7z3Czu6iFkIEoyPhG5/ShlnMoToUsPqaz+AbVx8hnn7vtAFNeXpUqr9E
vLWR/eIu9mxdNoPVlMNzzcp6YzlqiPqwqZ2Gc1MjxhDdKBm9rJlXT5xzjmg1d96pJ+znwAYSLPeA
VAOxtcxnqA+/mKWOLSNLSznXOVdRtZsrog1SxoceB+as8uadHzoPJklDyw9vIrIbBMyEU/bbnEit
lRxHy7cnQ8jMVRQS0oLe3bEBk/EhxsjkfVhUSRkhrW/u2XyR10qGHZWPXOyLj7MybU8TUUqtPFb2
ENTAVvS4uVlCNLyb34FTiaKO2K0IGG5/tqqzanRb57ymSJSEOJr1RxmLx1HRkX1fTeMO8jcRhsEQ
8gj42hoFUFZIGjrCiVdm2lVnb7NJBXJ07zecuwMEwyOzHeA16otFsBinDpxTqoxgl51IWfFJgBmb
xE59IaYrKm/WxrArJp61ZX1OyE0JrvXHQ9GnU/RqBg+16Q/HTtGwIwixVlJBaxtOBSHVax9+qnR9
kYOxpagh+P+gQZ3uRwfYGAD95tYS/vN63FMS08tclNyfGXc0CeVnTIHFHWpmqofN5uuNd7NeDk6Z
C4co5f37FumZREkrFWPXdlfmRNez3YPTj46LP+Lf0UQ6aNNedFv5bEcV3/HRnSWveO0aVR6+rZyl
Wi7np16mm0fF5xkHlASqoHMrvmbZ0nP1lfLeLEGRR9iQR+qqM+TZkMObCBIuh+JScwuogNYuaGle
XqTBCrhojVtoV5stIHdoZje34FYzwF3iWd7sdSY4plmiexw+VUZIZbArE9CRhgzlHcjsUNlGnswl
gg6shQguYLOUL0sbIdXQjM6BNwXYBW798bSzyAcZT5qfRWd9D2Mk0N7fF9gIkfdT6hfZRuAhKpY1
OElA8t1P1tqL6Uoix43uqpJZf9DHzIaZrOp8JVsLpW8yUzu/po39eJvY5kY11H8lFgKsw0MJt+Rk
JQsPtdhboElHJv6P4yP0mcamF9663ZO0dOLrmZxHINmG8NBcwLu/jfq7N99Mlv7wmZN5JTeo/fMZ
DP0M5RmL5QE9XVDLX1tUH/lD1SgXccTEPIv5a+3ZT7o9MS510n98bJ8AmaYoY76QK/HQBQVGTudT
y+v1GSWd4t5wNLPrCznk7yFlCB3MUyFA1aZtuNKIBvl5wDeUG7ewsi/3FJzV3bgXKBHEs01PwPmH
v4cqQZjQMTZJ9tQC77Vq0Hej8LilCFqjedRiQHRwQaGmc+kpkw+ot6CFKcM+as/H+o/UO6Ktv6fR
oHEB10Cm3SAElfnSouiYE5OFwjKOh6UnxwHLKVxZFGexaADlOfc7UEMuFNxH3c6t3hxnCA7zdDmd
EdbIxFGGffagOm4EFC4NBMXQJzPBwVnF3k4pWdXwPcOpndAIitn8dnlZao4mAirIhZ5G5T4cHP0C
WyCckfk09wJpialxdBuNNja4789KZBmQkYuZQSHc43tHsiz7VEmk2f7NZfD9gKyNO1EMxZnoeZ9Q
uItEZx9Pv8hMMB+Pnso8pMytenyqoM0lz6dzpdH0F93owsNNriX13FsdiYJ+Ryc6OIQpr2IjDFiY
Azm4edSDJclGmH1zVr3/UQL2RBOcJD65cY9rfBROb7VbuK9Pv4mn2qyHHpnAWmnW5cfPcHdjeCat
2xMRU6cC8yGUkLj89X1UfUk3a1WpAmefbzsVOj2XXZ8mJcp8LXMQ6umETvO5gE2Tbwu8dGyY916P
qV8B81t9SsZRMnAe2ogvtRRfeTMPy/KsmkoCHgq/jZFC5057ZHRXXXe+JjtQpLRdQTyUHOL95o7j
/a9cvl7CpSstVP0T63atPJLW0KmFbi2w4p8uQQANwyj6eckmYGVYFJwIhz/rIjGksRFvUUGTuG3f
RNtDxdh4Tj9IKTfdeUGIriGEFiSmC8ECnDYHk6qIDDH3K5Cz9d6Zkr9XIisQx8wED3QFzko8vZ9O
mKuJANEoP+nsTXAF7GZgAd+gRyaOikLrax7KuNc4YYxxtP+oeyAtFZUL7vwtXwP83zx9DIx2pkAO
SnvFY0jps44KT0Hk5FeCciZAWDcq1rvVO/gRBJ5+RNUNPIGP3W6W2xuwt47k3DSJYn3yAXaMd83Q
6/2dKxQPvdB47jlHBVS+A6iiqIO247N8bcmjKFwrrInoLRsqGBogPCnJBYAf74eNkOCeKqwM1E+7
62dHIpceT6gdxFjlTyMhnRPtwbAx9GZK2g670Un02ATj8SfwYyFEVa04PnajFsdRY/BbzBZdjLLo
yGIOwi3v1eN1z2djtrSdT26RWVbyDOHY+JOf2vHLsnDf/c6sjPOBeuqGS1Mm8kb2oyGZrmcJaFiW
9qYS1wtDRFiCfmzqOzhjQaqsXTARCn7o4SL+mYcsiKmS1MidCAdJxbT0DZUTdh0/f4/3aqpkPjAK
5WPIFFOZ3u80QHQMtFuY+Lx2AzRhWLt6nZvxmleJSLShC+Q/HIPVQ3/uAay1pV9tAz/mhTv9ihxK
88iUj/UtG2CjqVYIIG98w9xlxEZIiJVRWazBHTFcr7/QoJrzaXoeXmVlzL7AnsM9q7g+GxPX+JE3
ERf2A6mwQhd1aPKuzbxSJ0S3/0nwEroZB6TPZ68DwLRsJkdeAqTSomKPryfDRoBn14xS4ERJvJw/
BrbVjuDFn5kMhIkosN5QJoQEQdcrqrCF4cbIJxDFVAH5zgg9BIiLcXuDhHUCFGXt05vpIoRDTbsV
KUT0yUbHYpARx3+UBpkKn/Q4G798PMF1Z3vned6mHktygW6OCye+hNV1MZyRtethuEc7iN4XG2yM
k8Ve5g5jiWhnlqrx+UmWPS6tzQ73b33bwmJYziiwm4+KljsEkvRBD7ISTNF2k5OT5xcNXy0H4h8A
2xU8mObU5oF6GB3/INTBhINvYJkY4I0GsHND8ryCIPN2ttmzGU9JCjj4qC+U/c20uSAyTPDSVwhA
/V9YB8dsFtW2ciaNS2HWg3OwK4HzQFtJQOm4hBpaX0YTfxEHMCYMQKJy2Qt30JiQtVcmokWDCy1O
klgh8MAWzYlSUz8jXGmSirfG+/ZbeLF4XDVfmNRSAnQ+chw9u72T5LKg+FMH0d/Wl3WIMrU4t/pq
KDtFQm9GxfG3G7+zQ68QMMCDFH7xodLqAojhIYdzgp1pcmWvy+jv0VNGxpldX31hf0oE2aFa2kpE
6TGmRmHKZT47jL8K7iwqlEI9ZQ9sA884duv3v8n5VPzBPg+rRTDibR32JoKttSX4yh4gY72BgQQl
TOvLccG0PMNtKYVb1rF9amDDwXl4bzBf+H8h23NY4ROYbVAZ5NWlSNJrpCwaONe4db02DCCnZ4m7
tmATQBmaxceApwtTmURSAo2WeyUXO9e5YCweC/V9e3oDCKJZCGKs1uZN/iNQaXCeIlwUOcI8lq0t
qGDQrh7A1/7sdwUs25Zb2i+jlNlHoyrae8GMuajznsxFw4EUgla2cUuO0c7VoEbeqrlCdkmks5WM
K66nnoIFZG68dK6g2j/bP5IRnWSAJOhwa5WgZFXun7BxWTu7tQ8W4GsIoOu9F86hDJm9dy0R4w9i
b58QA0pp4toI8C8EqRUeulpX8Vn7Vof5k0NheOOtrRIrJz7IYTxDypklhiYWG3J2pkoiZR6Dc6mR
8aoouIbAK8zEmEv6C2DOQYsw29raJ2fFAoN6RJEMn5NfLgiGyNa5Yziqro2cRjJlQln5aMT2WHb0
qFqG0sCIYnhRxoIcyp0MH8SUSCYe3vtbM+PUpGu/pAgFuCJl7RYU8Rc4FoQl+/g285cq+L72k2JT
LyD1n7kxwahHPHqllMvjh50PotbonE0usOJaojUR7z0fmdgH7rNdSiosMcuT1MuHDV98gAn0z3rP
eJ1BnBoeQZ3mlgdquULJ1KuCmO7KvzoNDRrKyuuip6Kftq7dQqqdHlb3fvLrhy2w11/R4gDLmPdV
D7zQx3a4Js57NMCtufqMcb5VN/zgw1Kaps76ARJRfjJDPntJPJ2wBu8HBKLAcCluuWDIzL9ryGTC
b32uOHcv7LZ8tl79HOdjcTIqLnoowfeThQeaw034iuXK1bYXoJMa2T7vt+5fK5cxYn8DanO3Edrr
RzdS2q9pYfYm/tW3CIGT8+iVHW0IzHUgr3glAofEPRoD7mL3kUxfGMI1WqDaR3OWq9nTo8ddalMB
TxzRvIC6gLl7PbT/zMb4W61oUW0GT6b0JHQqU+Fo6AVlOHTTWZfgs5j8zouFfyQUsfgpFrX4tx29
LNympOq4ljeztYTWQTdU9E1CCP+QyKaryghQqdXQAi0fB4XGAWQ6lO8nbTy1rVOrJle50lJ69SfE
Y3NsoVgkkW3ZOpM9H1EowH24E7gllyTALM1NxInCXQgsx3zmTJJi//Dc34YAvnVxDKHMwmmfPKDt
c4vr7Hu986dxPMM/5woS+a8CicXTBTYGb+enj9wAtxJNBWJgOBCSSXAfqKX8s3witq+UA7ZGb/En
CCoErlhFLbhasCugoQgngKKszsUy8lMJsY4qKj9XXZ7F3I8NWgn4x3cYGF3N6CfwfCS4PDROR1Ff
w/JZG3eEQ5CQo3dxt7qKXi81RBZajMr7ar6VHM537sy8y9fztQTGQB56wJEcc9rFuLNlvlArzWo8
5f9BWilucZoj4DMABoUkYdDpRh5r6EgzbRDqXcupMosRqJ398NH8E/aFDpLzpSkxxk2utENx4E0O
wQRT8X9DgvAEkz+AfREnrOYVRa3U+cDmYQNo6zeSK7N87fqcbCJkql/ekCOK7zjgQK207IbQ1j41
EANExgYn3FrJfWsNbE3/bRTMqv8Cw2aRuTnEx9I3qlR+Wq2BRl7H8j4mq8oo3BXsknqmPnAqjKXI
no5qHlHSwngEFNViqNHmhLdui5cM5KotavbmktHfqU6QBU9l+eLMkKpDvVzatDCwi8EfDD9vQkaO
O66QFXmfN0DtMrkrjNx0Q/6R8LY2QkNMjMOY1X7+eGF7cRMPgUReFTCLSaR1JPM46yJ3tVy4Bhhk
HqJWpCY2LfC222oiGDRT86cfcnDKLsHIdZjlNcZs4JFPW3lTGf+Gt7iJCuFjaSuyjdmzCEiW3OX5
kAUVgLyokUd+2754rH4IanhLTPMZkpsOiJSMJVqAuZAoEA4+6agKgH5U4DRY/X41DXS/BNIPiE0L
3UkPbPlMPAppap4v1WqmPeCzzOmoU2o/+1o6lWl5xJ/+f2GwCp58lhxBi/4SOwDT8cNp/su5HnIE
JEWyGH9o6qeF9k+M1JmRgP4wC7HHqqmlVSOUSaonZdYSWEBL/jfMo6DE+NYROpjoGzX0hQ72Xq8X
x0+3QaxtfXfdU4hNcUesf7jD7xzREL/k9TF19+5NpzZHJYLwCX5k0sCBuS8qnpGj+oclJGNVzMXi
r1dDVQ4Jl1bhaxWCCvqkSbT5OyRF8yMBjD2XxKVap1JdKA+Y+62Ld5ppaB57vrKRa3O7tQiaowgU
kNIZHH1e7RJTHM57SvKlqNzExkQvOhGQbquAZt9anTZHlT6Y6GZRtrD/wOQ9Agq1E0g2pEMscnKJ
CgFM7qGSP8lgMSilfsJkUW3/Dwf35NoP23iFlbVIRSxdDqaSjH7CfcUds4BjGFHjLpNZ8pIGNqGl
k8RD+X1AvdYo4M/aS8njyOS7XxVGtUdP08bRetbWXsdm1JbMIXUcX4Mv6xLzprZg3yXRX0ulaurV
a+rGhzMHOjpN95HPj/AIRmbfD0y0Uaw9OOQXYk8rGG7jw/noVf00GkbfyVOMRhDoPRFWpSTRO3RF
JLmMkNnVTQBxbhrgUfpT3nwKpMELbUVtiIarvyqzFQ2h4XP/CJsfNfi/DQq45DamZVQ6FXBgGNf2
miZGe8ZEro6GANsKgDBFRMqJLJnqbcs6ZS7JoBtYpS8yLm/oS9YxF7M7ylG8gPz6bOY2bhW2rURI
tYo/rzIDRdIuxoqilxMIkL1ZNuX7VqCHwcIwN2pAIJFjCq6PP2sSu5o5m2rVrNn4R1SR3opgFYHe
9rndVO3p3qwL5NLbnl09igVGrlEXGTuSXwSzEzEPfJ8WHFBjSdPq5qwPZssLwdk8364E77gP6Whp
2bUhwU85ymgURKYRvCIp16jIAz42uTPWIeXvaPsIsNP4F3WI3aTVt/jxMAuAfvtDGy798s6bemqw
U/F06dJHC03Rneh9Va51AweZFbgXp7CE2e1de1h02ToffoRVSHD9T55nnI6dbOnOou05hsEipsm2
dQERW5NKSuhK81g3G1kVEGIAKhd2sXOxwqGU/4a+9AJN/F6QamVtqJ9+4GNUAqNQhSRkjyp3zyDz
OXS5uNzVlGTunmUctTq5ul0SxDgK9Gn1MIoFoIApG4la8DkgAKYbcQYZiAySNGwEuKZwHPbQ/jAm
PfszlKJCe6XhrfhvTZ6Xg5zWTV5FXwAQjeesU4sw+/1mReBb/wC+KXm5wYxWhZdqrTuvvb0rsY3/
m9wTkMVQ9heeEVfwXvURiTOB2gZgnAICiXq7YtB3aoNcshrr/ByH07CQuIqU+aJ+dW2MztCZz79U
KtnM+GUIz9/wHeDtSlpfZCaEIcmODGJU9nMr/a65kqSpq2s2PejeK4pP8h+GFRS69D458wP1L5YE
y0+JczxZupo6wzM5w7bYW2PiuHTfuLiu7rU8jVSSg4xw5r0bnUnYq/7Ws+bAfqtwA2TF2Kp8L0Ny
7iVQCbJ+A5vcBeskqDP0ub3das28ci4E+J713+uJP4eiIpRY6pJoVhjSdOF9JiWTdibAEmL9702a
EbHmJoDlAlIspSwnW1Mha2EeEFNFctWKVfJjVeLviXSI6UrVY8rOIpJKY/fRTNFEIFJiwzwHDSEd
VNB9Mlfth/7Z1qQL7RpHv0Ns9eI7DlyRKoPRS4xxIQxM9V7bLkKVC+oxRBDEe0FA+KeiYsGIy3gI
Q5WrE3KL94vFTqNJk0Bz09R2xlilS8baq9z4XKRqPj+LgQbAYK/CKpQHQ9uG6YmbXgiPJFrxFy6w
ZomI0fggLDyKAtVZCPJgexfGWIuxZbp60ySwAg7JvqGlH06FnA8tTEBoWxgWWk6KdgOcP+OtSBEE
RCzs6cw4D7h4AFM2YJYLriiSjbla7yKMxpqtMET2xMUPp4iu3c3rVnKhHMS1mt03T5Ff/HMLa6S8
8K6faZzBGIWJjzXgPVB5RJXFzTiOD/s4q9bkdfxvHvvHwMxs9Un+xwRa/lp5/qatjSBr4I+54hi2
A4Q2mfAw6pZk8WowI+nZXhJ5Ov0DbY6S0zfCb2vPWDs5aYoEmAmOXT7gMt/WpRQu1MIW0WViWETB
MU4343uujXsC8YgCSfXtxPnxzwxCmW267oIPNw11cnrEBduwRlxoHYAeUiLDSVV2j3w13a2sXkiT
U1RVVKIKQS+fTeHFI2S8l42tzBW0Iq4vy8GPbfIt6zY1bLkHMauZxVO36xCk7mHbNPrTFStxNKJw
qQOaNtx4CMvBH7LicyRNOr26LYMLDXYl6w6VgD63EQ34RkbhUTjHxs0Sz2nT4s4lscwagMv4q4vl
Z7WTEoo7+Gl0JFJGKMCMt1rABgIoiuMrW4Rzh0wtCVZyljSVXbaEMAo+ejh+vA3ApwgHbEVcsQ8F
Adqibml7L/l8m/MDMC0grcQRiz56J97ZBGHAneCzpIAY5mPZO6oeMV6c1n1ECJYtiE9DPOnfSw6c
V/MpRh9E3VFjfdFBpQ/LFLgMkyEOp4pmMMVh9lAvJux6eQXY1qMfIOYgNsMsCI80kWoia3KV4huC
z6Xo75NZugBnHDcKvbgrW7sbEsO44QmleGuxUb6T/VPvEjrrIFKZenr1/K9WfwynplmCKn+oOA1k
yA7VXS5XmAPXwRM41mPnaTlgVlSYZ3q7HAslaiAg784/yoxbS72sOY26Ls9+sPtXfWKSAMnp6BJb
pznLgNloph/Ufh66UIkOJ3zSzefnFPe416ydsBuDY6s8A2PFKoSLXIyW67lCIvZi2Y831FDwMYLb
quvsS1Uz6d5qRfdcAaKYOTp8xzEpgORa334umwQFCsUOkTrLAX/Mtya4rAApQlVIEB5FtCWj8Pal
KwLd3OlBHl7yhA7NaIjqXgjxgyEQeF48zQ/V9WNdHz25m4GvzPdkmrXRfFfAsMPSLzExzhBAO9TZ
6j+jSoCMxos9j8HOGld9LCjk+jqbc/cQoRdLw82kug14bE3DgF9tOtgsfZXgLMew+s5UIU8BGNwq
uorIRT6lGwwBkaB7zTk141P/7XN9qrBbc2kp616WsfykS07I3nQXCuNMcwl3j8pyS2wvUlRF14N9
0CgRBRsHyV8yGmbwTLdYEf3B2rdLyuD3pfVcVhj8e6EtMIXL7IHK+H6hAcVtNIo1LuXH9gNGbZqJ
Ple6fYzfbtXR5iU2o+zUH0k1ckOTKbvltqJP2Mp2iaCl8NW84HwPVL16Jr12v8geuqkblEmPLviA
N90T7MiRFYCJt+ngYAiYLrW4SnhO0Ba3ecrG6dADsswsIwBZjOiFl8wZ8cwSviTcnimggqk76U4k
F1rK8Lxe28lWRVVVG0gtAh6TSESvITVo/YkvcuCnlB9ZcxCH4jFimP+tr39uNEY8XryoO0qQiMZ7
5oXuj5I9B3cH44/uQWdwZ05ogCYLzM4fTftNEyWs9i0edLBG8Fc1pAAJvdfA/KTdqqfLHGj4QmJF
8cuXpXpluO+v9J5rX5RoYpumQIaPE4uNydY23k/qphz9eWvAPrl9hAjh7T/QJKVh1Ciq9l8cwE8O
XsB2Iaw2vsIUHd1okr3au/eJub7AFZEWfP+oAietxwN+qvRGxrd9+gjZQKx75TH+OHyNlyicJ7An
zNpmQNKjvHGlGWiCpIlbLTuxtgkGXQgUde8Hq/+KgxGfZD39G1evtaolUEsonXn9ZQK/OewE59vG
90qEtEgd2i4jVi6DeMYD7lzXG1vHXk3rdkdRhJ8cJ94FVjo0zN+INXZeA6DRXr63wvMZttnVbwSm
7ywytsiMJ9yUkiB2t+PZDBilMhoI2WdXCWCMv/3HmQYAbqNw0AIFdBCwXXEJmXP2fwaVLZil376/
sdKtrAmAJQlspvsdSIAHANAYTM8mPHcFkXNVpbjHibhHy3pKYpexgQ5QhibngvvguT8p2F4d7AUN
5P0zRrJHGqYqmM6Ecen/x8njnPRH+rkM2HzvhndcJsedGGUqlSFiuKxDXlwnnt9vKS6MRlGKjf/B
aBOncnp72jVtxUBSatYG26qiEwpGYcvjCO+Lpu5OxVdZzhsd/RzVLMte55pDLenAAr+b4IdkEhNQ
4jVYjDyr8Vdm+nZ4Z1nktlZj1WZgWHv95A5jVQwsCG2ilC+29B29CWExO0vpGFq9QAOd3esmi5Vb
4v/WZBBTL0n9Rt05Y+h2OCx1YMLQ1xqEu/Wat1PaP8H6mte5R0h3isAINVva5XFFGZ3nX2xiL6vB
GLSeAETXU5rSsWRQxx+WHsTA2pkXkprw8SIFk12N/swJqQgS1LZccP1uSkFJ6uSMqkxbwZcUFKUj
EWy+AyG92pQOjz29ggmCdSOvuFCDipFRjeruqvjMgXUiS7nOxdXSdyuK0nGWgnizj+UDpHTeTXtj
WvYWZn42e4iIPpHs+7K0Ou9Aoj8oI8jAqC8UCnRIi9mmyVIEmHL++ZnDp+xo/2ZMiLdhwO4EGDgu
OTH6ViTAXDMQaiAh2nmVovbfDal5fOKFysLmjaob3KS3K90/GK4H8/f7lwK1sLS6ibN+32AMa4Wz
fbhyjL/PKGq6w/zQP316fFmDlUwntcMrTIFU0oZwh+k/TLlL+SugVrZPwdTw2vRPs8FJTeaoHJ8h
VAMnQACtE8ywZDsCcr4+SesZKxIlbS78T+XSJOkF7/JEQNZEHgBE6MMlLQZs2AWZfLu1CdxqbE0V
7Ca1YXv7Mc3cSMwqKiEyekiaVPmilEkFSbeIHy7s6Ja3Tiv5mT+5E6GGF4xqICrJ6hO1c0ZxD6aR
7nwXQr6lxUWeYbQ72FQRqEmkeec0aR5q3eNWnS7vtYAF6sOjIWwQ40ByUnRkhqT2MsBmUGLxEE5k
RpDVsLj/zp88C2z855SW7tazJA1SClAT6xBB30ezVToel4n4gvGkOybLH+D49N0QGdy2RBVG+jOn
Y2t8FBsAM8SpVQcClD5AQfR2PRHqnERFLfXfOUS5PhhiCnJ44ZhbytUJQUD2YuF/kyxpN9ktnI5c
INsSbWdPFRi+tlsRoPKV9stqieIwWhT3EI3nMYbp6JvQ6Bbz7gTcLNZWhg2RdniiCA8RGtj4Hetz
bDu7SjTSq2EKXxRGbJ31YT5T5eWUGs+gOKkvXbaPauLGit0gcAOkam7dfrDT2ZnJ2GvWSozHzemS
e6qu87hvPXMaqY0eafhU/BSy34IRxPbEbtNfFzyHIa8PVldg5v2EHHtKb7mXTaThIYPAaGzNdPqP
8cJ7ylZ5p/CGTzWbVfla8G66jpREvM/iL323kFygOvBwEbHCvUieAF/YeD+f1ow66OB6SIHCuyEb
gX7d1/JtjWHX1xEI9FIv7H4FHYfm+O0q0W6Iijh1tpx94Zf4Ilg2jI/VHTFi1OYeb4YNTps4ssVR
rc00C2P2Pr5gZEchW56GKI2Tzj+kvdBGoHeU2YYIRh3oZb8WC4cNPjbl+h8L7TZvhB/EYNFq615A
Y2BdvZtDVZq2w1iJKrE85ZvtYoS43bmoa7iDEnmqsf0xRAqQcIEI+dL8yjGMAFfVxc0PfEjFtve0
E4Ya1s3OrMmAJDjwioSVvCHcLWZR/2rST0ljBuaKqlTkdNoe2cSy8ccg6LD/fGevLxpR3zPbVGBY
lGlS8UmUZGcTidMBDHw2wWtjlwBvndVBI/f6Zfp4mZpbprml4nF44KCPs+jixIdUw6oECvL/Yz+f
p4F1tppuVBnXrSpe1w5MuqAinyFmZLhARSERD3oCxtWrXCJH2YrsvR6aPh8HM98951RDEDkQjbPv
F6YpAV7xczmdxpXJ2P+EdBgEGn2SiObW30+80aTNQlXrmIOLOumXJwxg8tLIr2EK1drfFbTjvKX1
ArY6rMNtXqo9AR9T71AGYUGhMvh1CrFCtoKli0rCEi0coSGuPtr8e1+wEOVsD3iZbheZnM0qtJZt
mn9ZHyBdzGA6EM5oqNbwDJ/tLDTEiEq4CtLCLiAUESGP5vjiVBH/7kWK/fFTxGYvXQ7kem06D01M
2jBRwOyw9gnxc9UYtluEk97uS7J6xrFQ+zhbUjcMQ0cMXmdPyJKdI94s84Sj/UHq3bcXI9iPonB4
zYwHr6k3lYKAcQGzAM/OMMnREoFa2rhoB8n9dVsy6JgvDc5FP3vfcNYdpRmQ0bclfa7KCwFMa2h2
aw3FALBLiBtl8iatRBl0VAUZTIxW8KwEOV5kWKm9Lrm4PmlXWbvY665feXtk4JrxbUyZ/DfWEeX7
s10/6z38QUzjdESoZUKjBGcQKNm0wg6QiPxq0Fb1sH5crM2k5nafJb2+a9yuFvJ54OoJNNn5AhWJ
ZX8Ie2sbAMv/A2QfjqBpfJ6OuyuAmzUOaANm1HrO+3XVkmUBfsGQLOsVkppIvf59jyHicbhlx3gr
I3RAlxPSSMpeQywGzTrdjmx9XsApdBVfK/KAG1fgYEs6LqnbjnxR+DPycSHo2j9BJ7NLqhfhPmzs
Em3FZrzETOJ+x5zpNvn/2mioRGcopWmZONmIRhEeIMOAAmsG8rWxE8GGeP1we9DyWcAWMTYnVJxq
QKFyTIcrVurHv6r1EtNdPI6bVLQqhR9TGSimj6wl3bycD4m+iUA2zedU7zeaAIkXnGciPEQnRctc
/QT3NOlzlvryVVohAVrz/5dgWyP9dE2NumDxkNEHmaIGDv8fI6jHpsS5eU2RJVBMFVy/Vboqrgvx
LK+8VeaE7WGVROfzLTx0n2UVW6wF39jjBjfhxkB5DhOHqtJDjZIp0IGdDQUs5J6E9yHD6wd6A5bB
OeHDY7WqJYy3c+V8sYDaMsr4k2ITf558f6rjQ/RX5NLxEDTCWhrZfOp00cOA21ookNZeGfJNYCky
UtyXaoVEKEf56seC+qBjjK1v3ejiBg1kqeOEMvccuR9ofm3X+ml+UA5Aqm/WJA1C8hWgkGdzcdAu
xkaUuyz+dye3ZdEwUYpRDVcJGZhui0/lcfr+Z471voCwBYa4z3QT9fEb78T9zpI7qVc04aS4554Q
nJn6wrKiXz9hhUXA+oVLjF77HvcPUuxYAzMjHudKluqhbMRABLQJRaM0LJG5lPhcyzAPRhbNLo7S
ZDIEnzaCcYREmQAu/CyUtJpNHiX3mhHuxQB4FC7tI+PaN4s2nx2tSTm51AeNRul4W1NPQyRZZuWF
JYfJDQQum7nYjm0zXTuV0fEUKotFmE5yM28T9PI8yjgA8ayMWypdAGmZT25ud1ZktoSGbK9IgGmV
z+amem2JdGW8QtInb4rNXkMOkTIhg1TcrOL2G5DR7Slav4ZBJ3sIHjVOeU+GDmJjxnKvfVv6Ue88
osLABphL1GE/0TQP8f2OT+/BAuOAUQE4rcacm93crUzWZYnVya4c4TUAvU+XVWHBR74JBjGgyaPM
0JeYAI1NHREuiXCO+JP84dLx5v5dk7aWIsNaIm79VDB+oJrsti61DrnISrMZiilxGTq5v7gqwjAd
ymUv+L3/hT3bsNymhWrPELsUBQS1tTvxQGl1WoRrJBOMqqVoPcTSQAVNJIPagHoQMKd1ffS0mmm6
edlzzVNc9EnBFY48lh1QLFN1NCEtFigfMw/jtZQU1SCEsrb1Kq08vUsQ8agFV2L3hYL6QmYyKc4e
1c4Gu/Bl+SNd9FP1JvBGigxOcWrRCdM9PyOojNKpbYjAEaFkhPNK1jeBmTr20aZRj2Fqd5Ca+Ev9
MlW1N9W+IoQh0n44Aarp2tOus99tl6CxWixecYNr35SXe7vjZ6r9hVUrECHPbu+aD79kI4twNk/Y
p1do6iRhOKzfg5/nMIRrwZPRSSFZhApZ5SalwDIbUTXIkYgJlyj7FNKWM8NdmuqRQPISyAbHY+SJ
8bq+5k9IdmIPoN8sP4t8uhsNffDjiSCMYPLC7IT6mhrsUDnAcUscnlIX6J8hAd9o46Aeu3ZI5d0B
WxSNouViqXq9ca0C6ww7H/tuUAD7lsfChkYtYIfxSWZs0Wa7ny7COGMDlYvPiLLQ8dkZPjz9k1Op
YWiEtTBPm7Kd8YHnBEHmNnOf5Ttj/rtNBl7ybXCfivW43ojvNwkwPEzWbpSeRzHkLAA7Dx98mpke
CfqxU3j7SbWOEDxoF/vMwcoHaTb65Dx+lWHTHrnRmLXGDsLjyF20Y9s3t4joYlRm/t25q6lUxeev
Wy/iazVQyUIuUenEIjZTGF1avx//UyjlHHDXggU89kB2Pn0rGbdTs4gFIpfFf1wJ5r1I4nK4m77A
cvQfqpv4AykoO6KxUcfOU0+/Gio9Ri70Os+QVbYyhI6oTQQZtAfYOQdZS5fu6dF6NoVsxlQmRmng
q0j9heAUg0r05D18kDBHETaZQHY/sJlmFkOn1n6F1y9AQDW5V3xFX/kjL/Q6rsu2XZFH8+Glfg5I
M3eH9pPTyNjSYGgP7BufTr0q67Mq/s4StOCO9VM3IJYQvi3ht7iB/qZQwy6pchHKvnYg5uEe0b5j
susmO7oyii19cG6Ozktzf1MBRFWW7O92JzeAecMdE2bEhWYYSPBA69xe0YawPxy4RNtEnoKi+NRt
5HcNr8+34KTTK0ZAWzc9nOcC87wsovbduqwQbDufpnbJ04fnSManwCYvoSg3+by9Ayxw+A/2Ftos
GaEhtTuJSq9rsSZM3LgFeWccyGSLnTtfRCRUFMAiH6eLMZYncNxGU6XBR78UGy/M6SfjdrpMJa9u
aOZigNA+tLP2hgjwL6dgLdP8Thdq/GVPyR3H9KtCmVWUUM59cYgnJOeMjV86cJEmTwlR4SlIrQJu
vSw9M2uhVp1xaeXTU2s2EF5pbfGWu9XidoJHrxKjYlCqkgEhXZCjjbCIKyRib9sXiXd83rIZLS2k
2QgCWTQeWFmId1a9romCLFpo11Gr8prK6gt8XEa81yJimzAYCSMMaZji/cqzelkJzGVSsTgaaSAD
D4Q0bKLIGOF8u5wQ1gi/AP8cQuS7ul7pfT1CLGp+Z/bDKKAh2gkUt+eEiUiqfczLxqxL3m7pOrN9
/q1Ohe5KfI0uA9yz5j//x2W6rS9oJ3tlWoHU6XVGWnx8koASxjrgnTwRRV3cUXrvgTxEwcI2tNik
LjUix0f1D5LSR/lG8eO7hJTor9GOUG46A2auqcUaV8Hlahc+WeGxDi7oZExxSjED8LIbhoLpQ1/E
zF6zsFEfZlX1QvupyAZaHWHqaAOKRBPHnWPtBr87oUCdRI8J5jzetaTZD9M0lS491+ywGwIC3MHs
LckMb0Wv88+CHBlAv9l5Z2+1Z+0hk3aJrBI9fRkXAdr+zwYM8tQc0kxeerufdNEs9/qDXPiKXAPl
n7vuxgFyrCd/ZOmspDNYXVv3iWKXWGcQy++TbcmpUBdQepSN7F8SJ2u43IR6lRGrXn0rrFt+74zB
KSUkpv+fWqicqrDQYoUWhboR5NJtHpewq3HjCTgtFUboRPtMsF4OSz10Yju2hJs38GjcwR2D5YvF
ZTf7jgce/V5tz4fXoe+IqulBWqkjBH5cBFlifrUTuxHy7QBnFwJal+FvL3ZBHW4QnYuifCLeRlOs
24AMD3dklgGc22zj/7+UJXR4L4lBX54vSEmm8KeH9Hll+KcJv6Ez2ui1kyS/vMp85+qAz5ghPtN1
+0fg0AfQM30o0TET2PP3aHlNBd1mfYwbeNQMyDoSyetydR65hrLB0bmWTc10c8UOVneoOGqsIJrt
KpS1chSPN4kGK97Ak/3ShRqyOW+i+WJH8yLO6No4dx8IrZbDthgM5ZY6DLdHqstEHt2mAWDi2Ykk
sa+e+YvNFvFw3puyHHG6UNIDxQ6D23otsBtoOe4iz4K33aoscVyUnFg2ajN+GoKWQv/kh5vU+rIw
ZIaKm05/oDZsDI5o737aD1RzzfkTf3jx+vvcDIjB+ZqUIFHRQ+d5I+rPbVPsKdh/3FO1CtzgbwrM
ekw4P3eCjop53BwH5rzZe2ZnOY/NshyMwAW8qajX+vbjuNC5E0d11jnr5mc48Qd0ADpcbI0EgiBW
1/zKg7E1cra3zCZuBb2y5vlrabJp0aRFkHSRupFHYUwSfpAzGOrZ+wIaKdtBSiYmn+RCA/TGXTWc
j/nu9TyrDbVEqj8TKU9M0l/vt8yC2xnn2aXJwWMduFnD4W/AE95z0ofp1I5UizTo3rNTV4sEf97C
pmdPmgnyCjKEfLMDjLKWDG6TGV/2qxg7/HGd8R71uYQfjPcAwfCPvaO5CSVG1MeXarucNnlF7aNY
6o1ZXsNGiPHNCp9oiaiDTgrUi+eWrXSOWSC1ww1PqW9njgR/+KRcDkwG1+c3H5IztCqiQ1hH2I8o
2aU+bYlWKdjbrQIF5+p/wUVZvxox6zmqL0lOPZUOiQveWXEhLmNvtcAlCGUBPxPTBjZtCvN7QU1X
ebda5xibnKJbTIJaHfh2pd7Ekt6L7qWncd3IzLKKPkmNhBkY/1FTw0XvYXDMeEGpm5T8+Oi6ih2I
CgLpVSJNSsbtev089OBJMr0Uia7plinDeheC+mWGe0SNzlh2q3qZsNcA9qpyifdbjKLvpEWLrw2e
8ZiD3TVykp1vtXlGj5S0B5KQHKTHMMn4fsfaxmSGNdHr4D0xxked8vFdTPAMn84+yjxBbyQ/8MnO
/bovUVqIlb8V2hyxjkXkCAGoMC8N88XDGEyj4C8ue2hL8Eve0fmIeOyDWN9wYqOs3Illh4EkL2/G
rRhUoopwh+uR7qLDWioTMwRcEQOMUpAIaxZxiO2FSW6Lwa5nhIbirO6DAeaoUYpKa3N2qcjksa7v
oncA5/YP72rSa1QeDeeG5DjyzyvCc9fPe2TFqCWHcRe8UMX/OgO+fpTa5uIayoM2GJaiaVikcsLJ
XkbRVUJEDIBTJf57lF7waeAzkFRLS9Z215Tu0IsNdef30D/XEE8XuFz0TA2WjVUx7ESkAtPmj/Ag
pSSBZBtzoqPsXQ3GfOGSl7LUnYK2tBUVK8EOu1niR/p/fxSkFA9hHK279q/MISv4bxX8gapB/wp5
nm4pJChQ1ctFVtdy7dtM2kAEb9eHegltcmcbAashdJ/urlJa2DCW/cDtTbkDy6LRsvHpifi/AgRX
fHZZ9wGFJsfep7xVYyXgCvb8QFY74ybrM0fRHrf7sdX6v4FvQrkPu+RbikZdvcCjnh36LnpAcjGL
9j2EqWLHtqIBjt4No9F3DXaYyBVGgzkSNqqKN8k+tNoTLo7jF4YEYIp06b6T33XiUhMmnr2UosRq
yQlmI8IOfRbhwJWY2BL3nRbrGvfM5oxcj0JaCs6aP6nAf5J4mKmvQrs8iNasUqTlFx93jnK0saZr
hafIyeN+qvZ5AWAr+fFzrqhtR7TSbT8d1sNyKiWv48iH24ZQ2Xq+kKDVPw/MsPGGcU8lSYwTa8cD
SbtQBBFZYxYbxT3h8ULH8jjtrsuXQR36ZSiRzn6RZj+eezjfxQDPDa91i7OEU83c/D+vsJqiK2vr
bXlg5A1hPT55j3j1kI2gcfSY4fm9oLZjcyFWpc7vDxvf+nXBt1+dumCs98lHOy0Ve/rCf9cV7VgH
UroKjq9BBwMLukdE+I8EnlvMe70t490PZbfLUuYspAl0XPj5HuZSMFkeGQOXOj1CMlmhfCW54/JJ
35KODw4hiOOYUcPpZ1VL2oEdzRQxv5tT1qllV3xisiQ6qYXL25Jrl4wCPEYyX7iauG+uBM08rT+B
q0784IejDcHVfYAnQmhRk1Zr4eU3JNW7x/oee0lHV6PhajSFVRzUluY69SLSnlpc5v84j9t20QGX
jhCwKBjb6CS9R4VcpLT8I6Drsw0OD9jqjTde77hwDC6a7k1OD+xXJvvCHT8mQTL6OkxyG6ERM/Sg
HkbcpIFSM67igOJQom7VKieOEpbaqXeUEWXmlxF7DjvgEPD6/+MRqU968CYIW26cOAU5DFCeAdQs
HvjpvUBLOj3lxZAlwnNIHG0BzbnAxvcYfE5xL4AKWlnPq5Rg/F51YIfnjBsD4Wp6mZa8GNHCEUQv
hdUcJiNdvOOGKIQBhuDQt9YdpYbh6tIGaIMP0NfFw8MzLKTjO3ULqXjztmAi0qNctdKdpD3fE8oi
/8MAJ1kAVFp8bak0IaQ980uDKZgGlN7wk/WO+G8vwfpUvEGd3MCy4WsNrQA2g0LoFX+hWmPkwtZe
ftsANG5n2bVG180sOO+61wK2uOuj455u+r8yOhyZvcE217UHs0S6r4CUiywV1f2oC9ItqGHsyvTH
9p+/NQuk0otSv5IXkUkwGICXra8vPfJdtLPCqSO9zWMhhC3ePEQHPy58RUDMU4stFuQ56nOs9ek2
XyqT7QF5Htedx83Ts+pnVx/lBNwGZz7C6TdP31RFKjgvqCOemnrIMdqlufCa2dB2gggBrrPeksXL
+kHFr+YGWMrTxTSqb7ZHVkIM62wcvIBV1rUbiWay6z0kX1n+9cqB4GXnzPfshHeLkJ5rMdM7tEDu
QacrIxlkoofUllj8kE39IL2eGV8qs0atXBeyUPfer8/xDMASc0wZQjLhsZXM9lAxjwIcCktcMAHW
tcQ7+p+8UceXG2eD05+NeZDYJMpzhXlrhdthSwaT4VuasxnCLYST+6fyiT3bAe/dgzpM3Reitq4H
biVdGBfLNDVT97TfjEp8t8ishYP7EnpdZbrYX7Yhw8/TrTPn0Sw7odnCrvyHUW7mm5b1bbA/nmjd
tsl09QMxu6g+j5kmeDbVDlhx/aJWCQ9haTtSsvFTFKUXkL8DFYn9sJ+ja0IcA927ZmPDsNguafOA
UQFhG1SHdommaB8pqBKp9gUoKTO5YM1ImW/RInckC63s9uyDwU6NYnSa/RL5FwcpwXb+e8ql4XdY
glAtw6bz+sZcwuoxOhCA4Zwns8OjKNepWhB7iHNuwL/FIUmaJB4VYsw2/K5hqhl1WkCAJCfVUucU
G1R2woBXBOLDGPGeFjagISBt7HpaS6t+preqXQ59Jyf6Itu4foNekeOTC7dN6Y1g4vKGVxylzP0E
1+qynEgzbgIpUpW52VWols3kh9qhUvUFa79DzKH+OF2iGVjI4AfNoZtUYBwN5aeZUgVQzd08V6HE
AwoTUHlq9SNldbsa1xTdJWKU4KEGwQF4cOpMNi4jvbmRVGKPscf4nNX0eTcyJxCwopQv57n7jiD+
WROT+AK2rXwV6wmzUXIKYfog/NBsQIKvaoMB1dqSILMNAkpSY5DhFjfnpboXS57bafm0QaysVWsZ
J0ZjCvQcMUSSPxBgzF7V83Hsp5ZI/HvAC3DAm7Wo7bjT2IzuO4/G5KMRKJzLPP55DmSVNPGFZOCR
TaqAjaAPbgUAx5lfrFrIqlqV7u65f4mAuwqjkxqRgj2UH0pEH7H1qvPUTRoXhD46sCHjAsdLoECP
ZcYTK9pxhGk4MPhIkog02Glgr8BAnqT63zr/IoChd2aVaL7YMOvwYUDpsF7kyv55coECbR31adZA
UYP2Sitye0l3+loXfZx8L2mI3PmUwY6YLWQkx6V0eKwseaWftOcTFkBkG4CM+VGSediCzfzVgheQ
RF5n1A4EvtYFHti7ek513k0xDgaPkfK1frlkvYtxC3eKRsDjppwq++ZpRuQrWZbftTvSjXdG5eQW
A5ZzjKaceDqpynL5jAwkhnn+xSKCHIeagS6zZ8XL8yJdiLJoe0+H6qxCd70IVOzaplJnoGuAXjGU
fxJPsoU1rqGT1ikzwZVyguYEYvqOl6swBQIZWeP8BDAhZsm2o2llk9WA+tgQW38SzOY21HUMyFqF
u91fuftLZPpGGh9AdgZXg3x12doEoluamcwCqmrcpMvPVRhXW7ACnQ/wr1Tm/0VWLgb3MEcN3nWp
20Sx87QkbJ1qX65+uFP/Zks3prL0MSgm1c2UAgqnJ5nczR3av5+REhGROfszNVB+q3x0dAViO4jB
ShUIPa73poB/vP2qaEDqJVv65vR/JolcoVQKrBj5QqNSXLBimlmbwCgoBmPauG/o+GCLUSTWm3AF
n3Jh6EQtwBnYPDoo29byM4ttaDMphFPfMCUp6zyKQ4yp712dEBc3CpxskjokYCBMS2GKYwfz6bh+
1u94GBJrXfHmWUB1sPAV0kYuePJVQaTzqM7Lm3VG6TcRqSKSMX68DBqbReEw8QtM5R1Y0sJvZGaE
HCvs2Af1SnGO4Q4LoudJhLJFH8vjIax7ltr065/NF7SSJYN+k3ls6mcTuJC49S2tIT18eFlUnvXq
jhkZnCmRijGO2WgyKqdNHK/bZmyDiPi0EH1n0tURmn58zpsgVJMRQpDP1cgP2rROYfQoHYnB890q
ebZ8b3HE9/icI8PooGdRNYSn5VK5IDNvgCVdE7w05k8sZhQc4bJjYLY2wyKpZ9CpEHDHBROT3MPa
3eppx93mdee6sJ9sBprz77D+E+kjvy7Vp7VhuOBg5t6GU2U/Bv68EPOYJy4+1/mcIbRTuPT1i3Uu
fhU1+P9v9L2LS7SCNCyhtVrJ3C/uqFKST6iZtdlJjGRiFCypNvuxdmWFMdQOMbMEujQFiXHEoEdc
nzcZI5s39aHB1ZjKBBJgcv4dbbbtGvOxjfcsISgVQX/q7ga6P1tOVvfZ0vajp0DW0IZ91VQiXZIM
MAfNJsIS846lH3EORGWKGIxhIefs9+Tmav/KkXwDeh3VNzksoN1TOBBp2EyvQc6mrB/dHWzNRr7m
QRGNhcM4dFxIwHdWoGMB5EV+unp8dO71tlQwLBDRa8gR52gUwhUQ1czwTho1RbUVTGQ5Lsx+bYjR
h4HwkEyC9P7L4aV/9zz44VQSXGSNWwd6T7WH8/LSW6gBPgqsZqO0giqF5PP8ag88JndCeyTBz+CM
3YgHgI0DwboR8oZmiDtZNBYxcxp+8Q9ccZkKDMpHfCzq1gL6cVDkMNj0dUH/zDU0w7tPg114KNeq
qjUrV+pePLv+BXf8dAtdz2o3H5x4PM5nnD/d4KE6XRKaHtopgXzBgAiht9pBBb6R/uYpzd/bnvxx
GWBPBE48NkscJPqKzbjniFp1ZvYEbESyqBgAD96UabXU0tonrShrmlCX4EeS8tuQMsQ4lAUWdbd8
vP0XWSjf8IJi6VWz/Fm6cDCyFz5PdVNG9AG6Mz/wyPTEL2Eqe5gCc8lI3UbIyIKbiVXNk8cdYRMV
4FZfw2/0gK+CF9rfCdliZ4kN/b4KivGExxqFeJO+kGWATFkAygWgDBKSvgwlnfi3qWyvB/oGaHyc
W7Y8axg/58pi+GXGgTRM6L627QNVppAcfbemxhCqFdmczGONqPcbTsxV2HmS1ZuuIB086vIb0WDM
t4/6EdYhFi1/TPhVM9rzPwoWwAerxBEML9au8DS9G/1JkkqpoyZYtzJZyZiZMl8em7R2qGs05HyP
qbCrlx4KABE3VxkMp8v9GQHJp0JozXJkhL9/ZCtfYzPs2SdIgxqdfGzPcLTHy2vQyut7WvXqLYno
GI0GcdU0xEHaQSN1clfZrDcNRhZ9HZbj3C/SiUN0ept2FrhCKKKRPJ4ItH4RDVQmIKondtD3dmfc
hKALwYZK4T9Cyf66l/vgVLDm+F18WQK831rNxygv8MHu+zf60mPrfZlMDu/e2QPmCMnCQypO317V
J8C7tmQIwYNRipHB7dWcqecSw5cxFVlnoTStf5HhSLL/TrFvVU85pd510GQvuGYtlhUPFZqTDPEY
LayzHBnWMHvujoRy6E+ubHZblTbSpIPOmOg9cl8UTOhAAjBoor69kMHLqFAnFSslIpN0tO+5dWTB
YXxEjrsa/z1KqfaVdVhplc9f1fKaM+xFDU++mY888sXAYIUI0aYTspUuA2o7Jm9NmD1WpPnzCrMG
GnU6SI/DmrR4BeLW0mJJQOGdoHToVq1CER8Sr7q3DlduBHv4Yg5ZeVHszcO7l3c3VoWuAYyaD/sV
XDIQx21hnJVuzJl99CYEgQgjWCEaidFI5ZRTu9Yx+92TBG+syQHFPfsQGbdjX+IJhFg/08nWzKId
PAE4PPC/5gkdsX/F5qSQhSfiSgsQI8nIlPlfo5BJm8Nn9cIkRLNG7Svc5305gpleK8UZQhCBzFv5
/SCMV8MgccqD83r1Y9cU/Kmx5a1GOhER4P6Fq132aX0hYCfdy56AJTNSkCWuRDF2SjDdY6TGVe6u
IWKaJnAQuKA8lxBvAsQjgLPsxpVP/0sqTtI4F0Npajjnya/oKzK3+P1bhSdaNWhsShNIloNcJ0o1
kSmgfCH6tzTJL2w3c9lJ3JHdnvFlGDd6nW/Da0R612BktpkCr7fnr4uL9fO3KA4TcYYFgh1pf4Ht
jMroAPaPktv1mRci9gDgeK735Ieh+F1+P7uEj8e6Oh6zZdrcM5OJtSwxkrTc/iU7Lfon0h7pUayC
VAcYGrK/47WgTNSPah9AUdipCgffJJlEndeTFbgCsdkDiCY+6w9Sy0IdATTqhxW74yW/vc1O3u19
wqTzkIM9uP9nM2iOvY1MQGiPcI+NotIgZlfr9wJ7Nbw//WvDnkzKi/npU7jPioZNPnjC6T64DV1K
QTH3wlFSJBl8hiNksCBaqloeMvVclAJ900JpGF7Fr9yAI0MSG6ot6t/91ahuoeVvPntgvCfgSTLD
oz3SU7Bm8XXwLs3MpMZ/cmoKu2HBzq6gLsv8V4Lo6nAJGcrz7yeloAchCM1k2eBKu/5WZkIFzFpd
lLt7Sa4AzmGUlH12+W+Si/6fyq4jXexpXaDARkSv86b3x2z2qyErvmaOS7JF20VxjeDH0mtSpX5r
pNnroPKZSwerdeejS+PE382ixesMwVgxEolOGznOI94jBa1qEHVnE26EYTlesekerNcMvNlthcfL
whZwW1vOTUvfYWQGIYnRChnG6kmKmFwMtF54/9mBgPiR3DuHt/CNLG92EHUnUSxR8PNZ6u4GIHwz
FE6GpBkoDEQFV7ElAw49DNBgc1wM2qV4W9V3OnR7Caj6WdaQYjLKY0lBYcIDX5eRJmIj3bWJKyWF
blO0CtavWnSE/m3Evwt90k9w7UYbI8B5+XoP8ix5ne1Tm/M5vzCIy2wJooyh1EmsIzdt0D9dqezg
Q82RsKIDuo9Y7E8xmdyGu3ZztRKL30LxhnJpLjXLSnCDmkrkLmJlwdx3ISq5ZTHx1P8udMouF38g
T0gB1pD9l8qgogt+Awd8HZQ5ugMbZrdpej0WRkVtGOaiR7+dtz7tw5PGHFbpABBOWSaXixiMCqpq
jt6b3UzJwCroTjs+6EENjItH969lMVOP1JQE9DCjB9zwN8ubAAFlpaBBl4obnaRCCAag7V7wXx8w
SfAJRtojK+3Rby0cHsg5jUuRN243+c8I6iv9CKLT5q8GCXCHNcHr96D6Ulrc2HVvVxvFjgd/5NHY
q/HLvwgqPhcuzyxBgxHghOyO0tPH0qQD/UF3+7/YBs6RaUAKc3OUt5B/SeJ6kOLCqR7Hn803+BnB
tlo468hLHty5i4CMut5KYbu73Tu9BdzTle3BF5TDpWtvxymLgSiGO7AurDWQ8sGwi0byOtB4ygs3
q02GK9p5Uw21vU5ekJFLpLEjFv8KDgwcwJwzR5ZRRPAMTp1xes5AL5XZyzoCJecqa714XD/N76C7
LeeMvJ8Z9ipg3RJh6ez+KtIAXYtcWvrGLkHnmYbdoB8sXj42YTB0JEiBvbWaX8xsQAKmFGAYbP7H
9RnVbHS3KSazOj4QjCLjAD5ti+fQU6Q6YZo2J+/m7Yy3PovfsFW00VhzLRC3G2LpqgvyrwQgXtV9
DzsC/2apPqWD7Mr23oUGd5RA2hRV1DBLiWlBoP9Fwlq8Cih+P8wQaqld8PDCU7N6hsF72bfVeUHn
1IlUVWJ+NxawBUbX22r10m/wsz9RhS8ZYiil9fDOElx8+/tNSZqA18zHGyQFsvHi8E8fUvd8Dss5
93i2yPmhU576fDZ4M1KpBUGGZsywqmNZ0YcHOQfmb3fz+6UmyCTROrMyditqd8dbzxKOxDzyeiMB
5HY7luSd/hnE4/DjIPTqo7iiCHa0RSTbTfBAuSXWewsF315uq2pvJn6Bh6LURp3zYUjP0SmVCutr
IHJlLZrEDwdD2s+DA+uT1C2DboLEdO7cTNklIbuli+rm2scrAngAAlYpVSweMCzezfpvNq98SLGS
b+J0Z7/anTevdWcscBLL1gKPUkM5t1MxRsIjnj9inLzi3ktGd6np9nHZmzFTpUDdTPDXhcuDflPt
wDaoajHCTDNb7sIsSxDrGpwJ/niEKA1MTG8jcSj+NasNMNxWuwL4Bi/rtzQDiVp6Zr05JF2Uq1DC
F25gi7dnHH8Fs2skdsVv1gpDrnB7gLOGF7NcROry0Segu1pYwqIdKMnzZ3rXc+pyR3vS4WWdSsIG
FJH7M5coQ7wdW6vh5uojbeQ6+DQWFzxKKkRen0sQjfMnCOKVyFSpHiomYDAesIMI/RYgEDtNOo+W
+bvBHvgweyIHb13MAo4rX64TeOhVXgI7sZRE9WWdLPYHwVqW9kDDY95WQDT5jEW+fTyKsm2d2MpU
BXiKsXcszwhXWWSHtflgwA9RYfbcatNmEXo5x5jcMMt0UpdesNbJixr3FxN5kRYlk/iH55SqT4g/
WktuXO37Z1LOKqR++KOtmFO3Oz5unrfmNnevoLaNJrJYsuOfNeOtIl17BQSyd5AFFpwhwg1DSOpn
JmX9qMBap7I2D7FpqYOsAvK2OxuLscvRPtiCQHgKFR3myjCS56YYV68q/khoFvMKvGDWYwqLchRy
eWzuH3k//v28zcXNhnjXubcke0yGThUWEBTWbKU+SDeweXaU7HWDKetN8eXHFZEZz82hUXGpbArd
97OaztMcLT7QsrD3UGldVp3gWPxtff8ogDYYA53jW3NK71DClDX2LeMQMwTHwg16xbeXC9jzGnJi
NDrj5RpMu89XMadtSyOpxoZc74jM1IWP82bRpurUHsCDFoJw6oMvPYbDpS0ls+xmYv7ve8C98G+v
SV8k54NW3Ym/hJgh+c8Ffd+n5opHQ/qG/F6regoO/CNRKC6j07nFaQjgwStjhqdp7nPEj06jIrk5
mSgqJEmCgibfIS3EAFOoE6Cd+PnRzQ3bAYUdX7BVt6OKqXiQomEhcLqbf/ZxAwyV59btIyW4l9PA
z1kFQ2b4mvm64PDN75TKduQRgJSV1kXKMitGHwucJlzFZBNsC7PF7gXaQRKyNgK7K/AKKWyMKzuB
6RhyVBJoIB5k+eg5MP+mJCSdQxzcrrakUXJZu+Uodwf8BLSRAobhFVVmyDvOjJUrNBSVnZW34PVo
Kfen7lkPC1y+bea4xqKpHMjBtFvQEERReuziM+/O+ryABlZgvix4z10ipYw++W1HqsjsA0x3RfpS
x3SY7CctX9HVH2un7xj4Gz0jxmoeIAuwa9y7a/Be40jSfndBgvAPhFC8OX3zo42ThRdrpYXdhzeo
0eNr7ulhjKf0A9m76a92CSnxLoanw/llAw6GpXSGQUT9BqSEL/OIVv1YXIJ7LV3fkq/1JbKfpW7n
QOcDcSMWzYeohy95y9+ALgQ3erkXIvOUN1aoMG1Bc1iw3Kc1DQIfAFm2GD0i8oLHP5hq6rm35Qx0
3gxqiVLLfJ50W11l0l4B9JQNazB8eZhP3ar4Jqewl9qzoELMJ7Ysdbi77VUoxVv1XjF2Vmu4ln9C
rbvIqpT75aUUReV17ZMBH1/prqMQC2D8uIIqzZr/CGiV0h2odSP6L+TVmSyJQkVXvXGh0w8sT+7q
Bmx0tajaMZmO1LySvl4JM+moPWhHGFqQXj634qKkY0+IlnmMD5nxeMTah4D1vYSnlU5sNI47BA3J
8TAmL3fYlmckU0hfQ1RbluWLQYAQYaU1qQUwt0zGc24kx6SB1TKQDmMpixPpm1gRygXSG2G6lW3b
rbtVKKq0zmTPUBonGOZrLLWuvKZvIWznqQrZYWWLyGDPh6GpN2nepTWRhbwRRGc5WeilKYYDnHHA
tcLugIsg7usr+Rn9TvUEfzQ4Uw/81Fz/Bu+lJ3hsjO9PTAxP2Y6/5Bz5hO9WzqMTsYBb8Op+/C0i
lYkpUiyebkSl2i+mWo0bTbgnIMKUlVQVDMUZBi2+YzGILQl9ieFuQXTScuOHms4DVSth5vToGWKO
QhP1Tr74rrZQZ1XwqU1jAJK/f8Zq22uMhR0O709RKhbTUJIzOVFxPQmDJ13kCb6z6g8zZvUFt7hZ
I2a7PTDdSPceItJqo9kFdJ6xik4fJRLGbfBazlupvNgISI9FLM71EXFDUCm0HJnE+IEHon9ncYUS
gPEquVk6WHTtCM8KhoNl8Hc40pP8BZCoAiYKccwPD71JHNHw8LpiDaKqh3eBDs+iugmf0WT8VZiM
CwGXUtlZymGFWppLBVGUWk0rSs4uSha7fIGhkZdexfwcQD81qma32zKESTpTaNaIvyXpApBO1rMO
CWNFLOvwvb2bnV7rX6QAOblpILjWnKrNzq1qWw2kuSV9vr8/4ii7y7n9UGi+JJ0Lm+Tn+wUxbWz+
h1hXNNzY5QoF29ezVkLQxa2StLpCEQQ1rSMw4uhgJtcRNJ884C/Pk4GHrYs3ZFjzlw+Ccec4yAT5
LucZwbOaXKTsoSDlwYBJ3zLa3bqPYs0YwNCE2BnSrCqZZ+FNR7mKrVwEd9NiGFNY2/Z8FUTeG4kk
b/cL1SDItM3U9lEkvbmH8tyntnPrJ6QH3eHUiRX/A5J9wMuF+KdA1mYSZ17wkfbuWNHEaDOxpTCe
OFdwlDHwaWU+jA7i9gXTCf4A5KyWuwNmVIOWOzHwO1n/eYOyum2m9peju39/azf5HKOaYPBKBAze
tig1g5TFzEc5ZdmRcWTeWf9kMjONYnS7t2in82Yzjca0BmFIIhreeQv2S4fePL1uPfXZ8Mode+LZ
lDOuLk3EODJEUQBeOKTGkPX6Ng8NevC5B1qU9B8khOFuYkd9ItueW/ngOK4M+3YKVI8K5qmUiyyd
sNGl1Hi265/QzO8W6Sa7dtQFWNT6b8aHWP3dUP0o4IohCaJ3yhIuOVoKqrp65bQiRFmXmsdWdjH8
UKDhMZc81a83Yz9jcfXdZMvDV3rj97eDlRhny81kotm4H3JJnRjuC4EoJgGF/i3ovkTCKLPRXSqu
G2NSrdpZptNgWIyLRHh4chvt/WbUWNqCKNu4DT2waDYvnWugM54dV10dadqMFvcZ0IeFgQLEJuV9
UwSNt8D8KzcFRQ5FDC9AjmnoVNd2L3haryYCVJ0F2H8ksiOr/Jk6YrVDsr95aDM6ZxqsVVXw3rPB
uO9mPTlVjJlCnG79YJZhyL1DiA0vMFBo10Amy+Pit2JXMzxxnOzGbC8BHAMfZouDR2YE61Ocx4CW
lrcwPOWFoWQyeVHXYSTpq76oxS3mu7qQkLfsJVSmD3eSmeOGiSiPwWiAu+fklSX6nBDpPTbvqpeD
I2VopEVj7uKciAbSTza8bzkBgqXd8VBmfgG4g/JVJMpQ7jqMFKz0avTQ6BJBfEXNIaZm/RqVlXxV
m2rU7WZhqowW5Y8uVhWKQWrX5DbSKdff0Qm6SoeiHBdwOMaSXhmxmTMG8I4AjKKNZJA9RUZfVPCx
mNWEuOZonmtWSvdEg8ZtYZRmE8biC9y0fk/MdSehD9HXr+0+uxI5ecaJo9zOKZci5KdUzJDxRi6w
3k1n73hxGbrBziOMGSJSvpBUr4VbCK9gtXOm3y3OyzIcbhWIf5KuEl1NBSpqzBKBC4GYuGLYRl27
rwj1dwrWLRBl7RujyuKEN3zceRQ+tu3dO6f9f6vPpls6aazA8dcZ3bK772l/NpQ2SIlk1Q7MUKCi
PovhsM4kawXO5BElJM1I4dkbqL076Er3z/uWgITeHFxGEglOO7nCACBuLTu4ppuLKokT0uRngnn1
Bk7X7fjvxEHtfsa2DstWQlIZdzJTx0vvJpJD1bXrHWcFjq3ykaBXe03bnxCPIstM5v1+l5dQfkMJ
o34G2AfqFOJu3NiRn5r7Vpy8tHwj9gl5GrfD3ZqtnmJdeEd1o14AI0gUW84d1ndQ+aPwuFR5twXS
gnDeVFer3109LFREFRetGdQLbFrrwxZYL7D+UeCQPsrFlt3Z0wrGhBTh4MjAf9XU9D22Ioi4KG0U
BRFLTaNzOMFHikny7pJj28Wy8fS1xBAIVUEYnquQ/x9YhJkqfnVaccl9H2oBbNLm8xABvj+EotlL
5iQ2mcB2lrjC1+HMK9qD7fSYpkhGiJaDfWER5YmxvACGzQnDgg8VauqhPc08BrdrL3SjU1uXrQ9b
o4wanijYaTShVtOuFzSFW8Tc3CsvWFLtXvu04c8c67qulQ1q8E6L+HdkSY26dziVRfIEx4WOaQ3q
y7ZOkxAGCoEdP9JZpzg1M22UDijOFyK7Ja/FjLVZaRpZEd1zJbdQ6CGPsP6iqa22pDi1SfiDN9nX
QjHZy9LJwGamNBHYjxu8BRo5cVOWWjeoG6IEFjg8z77dhKqQ8E11XhBrfmmMrfCiG4VjhPPDMLNV
OthL4c8cz1pNvd+wsF3tx9l0mOkivn5ohXx0Q59SEhjKbynQTy0pClrJBpqkw0j4lKxTkcCY1Cpe
DQHWwp5YZi1LBVN0OKkW1qac/o9r6CHJfXNOOkpNmQAh7klRBq3FDG+a+o0TdGB1FwIKeRYq4D5H
fJ4uGo+i1xf9k7f4HutWHnt+1ICe1e75ihDSm8fzYKKUuXWyQP2Y6k3OQk17rPCArpmdsFk3kPQK
wbZJzQs+RCkT6XCm1DjySvM8b5PY39VKsJLdZGP7pgGoQUYa2MBUErZnYiwlscx+crD75Clqw0N6
mvlFtvK6J8VdZ1Iq4kYHL/a/uo8m/SOsPGtK8key3C7Hrr35mC857RycxZOhgnNVLwOR0Kz5HPNt
cn73ZHSwNQNkbDfntSV9PYYqbl+uBGaB3Lg6TNBJpM155PuX5iS3uTqnW8TUwEW+Jb3NQ1XyXqkn
AhHoUF0wTEBmwuLO5v3pQAhhUtKijzwhezrcqLqL009Mf8L3sMeA1li3W43R66M8UD7VG4d9ZXCa
GxtMuQs2ILm7nbWbUtSmWtiF2PNVClHpO+aI9B3UuUCE+unsGuyNepLemykNaOmaX7qH3/nKPfoC
YZ0eF6bVuBU7o7aectCBUXKOjaO1+I8NrHUEPcNUKvXnaG45Wv/RCffW25c4TNoUvtwlTI0J9DKy
qN+sB94jCz8w73FkMIC/xBt5jRLjca9odz4RkOOuZgaNfwjjZADtOY+GTVizhV9S2qOu+cb8UtHF
QLoekMcK5QfSOE1pv+rvnM2+Dlwd+a/vSeBGGBEnAMOJ2DEcU+XCAcns9+rRj9Vs+zBh8uO5AOtR
mAnSyT8NqaCkpCEs8tptke762IBJ9of2imdiwDPjhJZYd6zYtAdhGTAGsePaS1M8kdmxRqeKx+C3
lKY2vNeQZa3wk4R9p02pKod1L4fEBNpAGHtlne3Z9MUTf0zo4TiCj2GcBs1QAHlBL9hyxbt8GfEZ
hR1gmXGlQvewoobBZ+sawPjKy71ZajekM6ECZLmGvZsIb1X94GvJYv3xlD+/vN3QVLBNjprMC8cY
bPgdQ6EZVLVxhpGICmhQowp+NYIdx7NUrdClxzlExk/+oKBQwziYptIFv0lscAxWR3xjfnLx2lRB
Dry+XYFiQrJKnI4nIAtMiYsXS4O1IVfa0RyvFzBy6HSVrM3UnnGTfzV3NiDFnET/SL/3BKBz19Fx
6Ek43aLTnIpcYXTqs9FTI32AOZ/E/pMzvBC9nUEtqReKhnkaZEym9szjd1KzmlxQoyaEO1INoN0X
G//el4A8ymEd3v0tTOprseqsnD53Xo/pkaik8uSRpY5rRtsaZlU3xl94DDzoJnUantk3S0GMdS6C
y7IFAp9sa1UHBco6MI+XeKQfWXZVVA+btD16iE51KfXhIU1TXVrpuT2gaJ6qE//iPxSRUvGTbsY8
kDbKBaA3e35QuqwwLbH3zwURTJbWmo4BNOIEwRpTo7o6yt/fzODvG07w+APL1XPfqE20b0wWmUSc
A8lrqxmAvZkpQ4SPY52AIY9BSrsoGvJL+ztMbMWEFBVpUEzhftAVuCjmZ5zTbXKJR+YbkWBQVo6P
//XYmvJ741DSuIu2Bgt1DXxboHlrzvjNeOghkfEKmTEu8c+QOk00kphcodY/MGulk+8fkSV7mQr0
KqmlnffQwAQtI/B1nN52KJm3O4KcOqy4XrDVZ+l0P2XzyReJSVlciYhyCH49jqpiwrKJ2CBOF8CU
ISjOkRwdFemlbTKyXapIoaUvKwx23jK5AsiYOZfxV80vVjXRvVFSRHetRh48A0iIu9UKQJuqjg9A
w7JwmLipSiMLpWPVRxuMUyxBgvhANJ53VElzy3IhuJtL+dbYOPMOqPTEM5j3JaAdu2cErY8OaS3B
Ny7biaFzeI0G3HLHT6fWointGFH2liW+I6DF1k6HY7o3UnGfwyXqg3yICJv8zO9rFxOu6kpwiZQ0
sO+M1DXsciwQJH1wRmnSrjpJMrVyWhqg7wqRVlBlFd88dUDDKf8Yziv0NjuBpaGPxd1t0h4XjypX
A0oyd3iYl/puCcuqKu5Ii7Fvk0Ou4MIv55Lsttgvgm7EzoQ9hcX7H64ToLUAIfSZJwbUnhqmP5S+
hAq1nLDQSWoscRHnPJAOYg0H/J6fGQXR+gDtY8YI5snOat8LFHzpmYpWNleNw/fUQFlZ1IFxVeCh
pKonWbVUk7HKzT4Z+GEDMGbiOjHBc77E0np4AaXnZtg9WQNSXk/ljLFqajQqhdIwUbfjkhdvhBGE
NHrXZeXJy+ihXdA66D7GCMuqYbEkal+lR0W1/NP6JnUaxh5xAqu1RAicmA7vVr7vMZmcZTWLG0aH
Bzns6zwxQArh6w7dByS5Krf8gVwQ3wCqJY7SVzUdq67JBaze0k0i4KiYoBc1vdWSxtns++VT73Dd
9jOh9oTA2AWYeuEy/G8p/2a+sym2e24MG9IsvVIv6tCMG6GAlt9Sj7RUYOFM5PV2j7sh8Fg7v1rv
G8WIM/5Q6AbOAqEgaypL5myl5ZDtD1iJ+LbdFLmygwZdTbYia4E6FxBJrLp6/6T+4TGzd8XoGiOy
jdlnL99Wr2sc5E9Cw2FyMM46bstaKOXAhrl0XWu1JCSyPElo3sawMcLSIqXJT0FZpJ3Y8eMsrFDx
FA/kqOaiJzaVIGhdpwzPsSNWi+erCLfK4ekmPFtcOKmmfhmLo9vwHlidoEzer8/jKzkm0A32dKkL
CogH4mpsY96UnHcy4PJ9RszTDu9tejhoP1ZzN1JHeDTYeTMd/ZrK9/JprUo6hET7ToHrcL7ALpiO
PSeGXVhflcRU9x4uVfRgIi/gKCLtB43XF2M7ZI6iuh34DquUJalUyu5zvNVxS7lnwWV44SE5YxRz
c2wW8bDCwqF3jCa4C3xvcV4LWEl3NgLqTcxSLB8MIfU4SNc3jqdxTObKRV2wPQAAiulpSBpQ+j5k
jvTEmk8HaAvqUoG830thd/rZaajYqGb6xkb71IbJ9CZkgWT+5mxxcuanvHbaqLZUjNVe5rp6MC3p
WRn/cOvTj0qCSYSAii+CHR+6su4GWPlaVR6w2npy8Ph+1Xl3iIJ2ojMoZ0UdQEirO48RfhzDf7w2
EWZ0C4otx1lsMtBjBGpSg7d9t6rC431M1CzwOQF2n1Vqpz8Y9RVjFBBGrUp45qQxXuVBNPFQ0nbq
Wkf2RFmvvFtt5tZgy/V3UJFcKTzJFuqAiey1YRPOBgNsS2QJn/+EykLUUIvmYYdu5KEXQkxl1CGN
XCSRrLpRJSyWPlnj8Q294Yz3oHlSj+bCAO7YGlHmBY3RnvxBEORIj1IOUNeJLa30ROsLPo96YPlF
Y8hnwy1+nA+EUZu46y1YeORupC2vglOL/2kFVxjK58iBa9l2x4N6LMOkMfJQnDn4++n/Do3a7oju
FVkAu5Uq2IciTztawSmZLOHRkWMcHO51V188YjvIt2jCSXMLkZTQERttbvKjivneApWJabGGcGoD
a0NNrlTCl/EY3ZJDdHf3qwWMhIBmZnfPadCGv9cbBH9u0nEXTEokUgYVl85met9AyQ/vevB+3rWQ
w3os59e5mo26mf2tpe7NHsBoqRFSlO5NLikYo98YOz53EyLm/E0VQOg4X1E3yafwv6iqjtPhv2oC
ZKnS2zyOd5+iiC8a+sEfvoeYl+AImfrsHaEKWe1gwlpUYShYFiEUnRZkZOAv2YiEArBDk7TG3G1r
PtSXe/ijq83PrhilzsV8fjD9d8+EfkJiS8yOCqcT/6Gnebs2Yf7qBfSEE7useftjqub8qx89ItPa
0lyl1V59kMt5PNgp1ZpHRYS3INx3rp5eu0z7FwtStEnFIThOq/ZoYpYfV48HPJo6wqrekkE1a8ZS
/ojzbZoTSVqFfAqLoRkc/C7d3ruMGHzMDyM19QlusnO6MVcR3JMcZjrmdgwyrZmOeSBvgZWqG0EK
YQ0Bv6ItrV1OLOfK7e9odxN0jxJBqMrlfFVUpj7sKteKNZsb6sYrb2t7TO4FxpglXErKZeu3bewd
3Y9fWtVR8RXOM2yofAVg3adNEnfLB0NeIArQIQtQJi4HUJS6Sve0q4vwdj8TKrf98Q/Ci72B5VK4
J2sO8b1IG1QWZ+empUyHTAYh89WSEUazK894pNz4QfHPQa0ctfcooJIn9dSYfBhzkkX5ekyEykrm
M9bg60592NDu4GjvN2fcn3k/GHlaqPsQ1lvIM5o4AqKt1gjnzteS0cU2T3qpwNmTUYiz6y3uCtlY
/KevyVq3D4WJAutYW/Qg07UGcbVaXofpzMwcCeh3hlNsoCbEgnEKcqWtyWQWv3eggC3zWVs7QMrw
SQa1UA+1Av7uwWn7hfzEsEEBhpysoMfWBiwNbDjuTitOV8IKqXNgaOyTr914e2yxiNG5XIAxb8sC
mkrrLPkd9iAzjX/RQ/OZ+t9pjDirIUvlcA6w2MSH4YTMnVQxPDYwNShsGPEhkNhJx9hAAVrCZ429
RC8tBwCSpBlYRQ6mHd3CeD0oE8y6r12U1H4tqaU8xS/c+BaEC+HJ8EyVHQCh1GHfSPivPTCXVXcP
fpVcXKFUveXK/toPH1F+JwDgtRaJ42y2U9KJ1p6ghRvzp7HMw+IvLv0/sjaM8MyFkV6CSlKtVStw
DEcMECKcWCcahbHQdIYKCAi8+K92emBfn0Ds/v/JSpkQun2dMDXLYj6Qo8OIJSTPROFQLoTNpsXt
auGKbmmpoHeqcttZjNbb9Y+jza+/As4Bbf7HkyHnI30vaJP4Ct2yuBDsDv6xNrsxo16u+kWoik1l
NNSJV16g3LDPT40558DvjDjOr3i6aha6ChD48CWw5nKeqHq/0qBoHt2Q7MAOj2g/LiixncwvZaYY
xQb98g1qhwIQJwrX8a0jXLOSkBYb9V1m8VE8UYmgZ51acc3yTGOiPPZbIZ3gp7AtC9CeNgsIEvOJ
54wJAK0pAe8rFvCQPh4nQ6UVSf92FLoJN4A9+tQ1bmC8K708UUZ0dH+gvZYfpRC25pXB+qqInHxg
KVF1j2Fbjp5YtcUWO8NwZnUgOiKgtlwTp1r33sLD9dYSQwqSGdcljI1iVwo20ezV4UYVGN/wm5uM
U5otg4RJvlRhqjJ0kIHMG/GJ4LRBHYh5jNkVXmGdoU9qFd/mka9fxqbMbcKWlqoxRwlziTS5lFhG
+kBEnW0H+zxSQ8olRuHhErkdwvDvWjtHpeYBnEW2HJqQlt8ucH/R1kbFU1t2HTwskA0zEVNJKyr+
XFPhc213KmKF3S6bvAdm+J3P9ayZDbuhDxFksklsxaNQO+TrjFX59ncMnulgisDLpff5vjWNCFoQ
/i8hWY+g4LAeV4owPkARgSx9mjNVUIWIv61Fz9nHWCz0PJ3euXivBpIO9KqbAHLqT0Cw077cD7Kc
1/ofTtC4JGkpuWI+TcQbep4nDKfjWCDSG+ogbvQ/sWonTBBvsaFs2e7QE0dYBl59F5ORMg7b7PnA
ML4LRLa8DTWZ3E4n1ceRGV4nynHolUROHFR2FQjoBcSN/+o5fcliMn+/s0ICouD1XuUi9wYsccht
XDf4MlnxD3RBLgtdaRAt2++x21C1nuCqvBtdgK3Z3OGfbCMjmRrR12yxEyyenk3a2Tqrk42BcDhQ
mSLhixPYOAZjq4bvsU8aJk2HUv5lDTiu6ZPfWcWb04Rjpx1y0+ANY2mBTPik1qtttsxK69jKoH6/
iNO+xx+8T8BRMCxf4Otc8iW/V+r/mLwEpyqFPw+eTPcZ591D8OXotI2xpXz6C+RaQGHRRydMbOtW
K/72ox7QgCpGet5LvqxmAEjaGGJzB7pWB3XmjZiAngBKcyzNqu9pgpxWalSzlJV+A+cL0dBecFMG
cgdb4rtGJ27FPMsLNu5FvooTSjJsbKgQlnSFwbkH31HyVDUov1ryvBCQGy6NVk9HGdY0xkDtX8T8
HVNtanLeVUm8Xx++BuFr0G/stdfXx83g36hK04bQALGzr4YNZ0mvVblb8RYWUolvTwE0XYAdJiaR
SNbaZSiRMAmOxCOQby9f6xXuugsXaXjRQtCeNRmwL1m3/CNwBOB6lNAGDXegiLd9qzFiGBy8you9
RreKjs/tqC+oa+n+ML0ASE9kMdsCHNgwFTXPPc2cL3/DHJUdrzilE6t6zwPmuW7vtbOyV9Cm+ftF
Rxstxn+ZPoxw1rsQH0u/7SV/22C6tgzPJ05uLdgkITYFEVGNpAzwP2hZ6aWgSycN8CQZFiPsnxES
aZ2PJYFi7qaR0Ugk7DqA8Rw9jkDqNItRYtC24k/3NUgCNbYSh0Wv6Mq7wIQbW965RgYz0zU6CHQo
YEJ7FCvVGtwJv3ITzotIfSZi06Tz+Xv6lghuy/15jECgMia+auFIodkguspzZjoLBOk6EJ8GE/KS
E/VwTPKG5VVYhe3dHqTkT8v8wq9LVfKKK4tOKyveVJX5pZcw+stS6/p7YY669XSatVOp6bcXSK1g
VjPX9GxyIj1YN3wglpTdkRdBYFeKee4wwlAfwWV8KHEAnMHhgyD6O1rVwhXiy1PCDFuKAtsbHlH3
C3ohaVy3mnjhagxMTlw8ySXiUUyPvVuiwSUiqVxDAtAjrLaRZIqcKVE5k0YxoLN4AfkbJZQzF73c
iZO7aY0aXRKfnG0MUgNDjxehOkw7opHTyRQcFfZRnZR02O8SpezjQBB5SAOt9UPnQ7g1GMXR4eXY
u+0QDG5kqoA6bph4eq1dAghmODVZfsUqydhtLFFsL7IFr3yq16ciLeow96sPu5jpJlbdtE2D5o2T
6Wzfg82ri4W3U4clQNOJp6YsswazTzqTBtGhyAELNfy5E4bdUgDBPfYMHFHVP8dZLW8hh3+q59KL
vJU/uQLDWYfnUiWg8XXXXxOwnHQuwTN89pzfha2IDlFBYD2CiB0epxGH7+0yZGVUxFsV08DyyZ16
r7MFIpAw1yFMUjBQijQMgE58IzsGpmNQrGMuajuI+yk7aV+CGJtgmnCoXRUoiBPYutowJuRuXo+p
oQ8sHRKmRg7udV3aYmalxT7Ks/6/Lti/zNzTAv3FHWSxGA1quJJiBGKl0D7IZYmTlx8LS1NAnVV3
+LCocbHzfT3PuiEWWf1CmuNLosFWfXuxEjidyqAyu3TxqpTuhriqVec/1HBAL6olKpm4zh6mrZ4T
F1Dqlc1tjDUJswYW/eEw477AbE58YxkVwNcP10PQ1L+Zj83dri/jzQ06I8DgTLYM65a0xcmiJdLh
1VmVlRGp6FF08Adoz44c4N2wSHRS/m3PdPwKB0y3DQ9EUeZykwREOI+A35u+/1/mFulcCn/PDgV/
3cOtlXGd6awaLvYakmSIKkKLY+4XUvYiC9w8d6SPKXjdeTG906kbi9ezkinz/koOWQfFYu1VgYji
qmpBlEkoclBZS7GYMyYwy0ks+h9EgNC+VXGXW6TtbJCkS68WkGXEm6lBLL34lf4Og3kEXa7HAcL5
JCyEKzs32mYMxU8w5CndWzgBNDa0u1mTpgZY9H338ygmcVUBbqIUeVgGwSu5rMbZZCX4lbca/xo/
yVfaqZ6CfTA1jRZfFGogpHNsiQnZz3XFOG0WZGFbXSQ6Xpoc0wySN8e7CVcGi+fhQMBZ5Tea0H8B
D6yl7Ov9G+vx8lxsVpTiPUdNI6bJ0fTcmw1yhgVAsDV+AFNd05AZCu/KE/LPBRcckBkNII+bF6RX
uU0Hw8LxWVSmFZeDhjFi4SPKQ2wUVakGrLFsXZTJj0ORsFiUCI0/gM2YopZMPfnhuMQ7gIyhEmls
JBg+oHQ0WO4UPPYF412Ja/UpU6InSh3uqecvXThmS9VU/HhAjYQlXx8CCKcEGT1v46EOIzA1dtTD
6gOkI90mvi/pPG38bUM+VDWx5vR41FDZFvl0EAehrJom9QKcGapFq3eRvMxiPGAPEdJQCP64u3+9
8D6V30vyCZ5zIyLqxlVJx8jsEuIkF5kpYAE27L2rhPL5IrkjPb/4zLB54+Age3CtjTjcX4jkS5dI
XVCrU/1x2w4AisXc5zmKUfQ0L+rbbInqOpgg0P7zriCRMP8tpysqZhiT6iBFBiYcMdhfD5q4xpaG
6QcZunmhWzniPcB61GIOS1CSRJpAxYxNZI1fAyfoHGTpErLGMtmLf5vFiHf3a6MTNkQSTx5PJvZ5
d+V2Rsx8j4pbhC3fBOacFOr6WJ2Q7lZkDW8kfoIYp2Sb8qlr3s/Uvfgz4pAQaFPl8quH4B4faJsd
WELPhtcvfApds/JdsMapzmbaGqXHEbvqPJXcgiQDqpQfvkg5CGlPthQho0I7EnsGwI6tflGG+al7
3Z/RRvikEgQUbWFFYI6FBVVN/UY9GSs0q2YyXxVKNJNsgpeQ1AqUbxhWQdnCpJLhQpD+wdx4Lbea
xXn5Vm6bPL7BMdZG0YIXFdlshJ0J116K8C5YRMIOwXCFd7N/EkXRxKJqTnQxaKlxuyTyDGK2qnzm
n80010Fg1BnkeTWn5m/WcVipn4rEN+EDZ8FbvTCPe3WY/1NyaEO7eZHV0WUu6j1n2MsafIWEsKKZ
BPKJe7mQL0wdgZIWztBtfjH5zKHqK5MX1fDVJ8cNxwHNtq97VigXCZGKL6Dw1gI31kKVkPWnxYXX
eqZDwVRSqxhl9mczzPOQaF+Qh7CwSntXqiMU8Rw9KroteZkA1ZpTSXGfbmnb3NdfhSaW1jyaiIhP
3Q1AYdBzyT4rhdXSNknIHZrq9WhOo+UWZYnY6JVBuUz1E3zI8jLbxYojgE+tcAiFbGqipR8tSJtC
2c2LQvcZ3qjtIMogGD4EogA12tbAf7N4W787WPu9QvEo0Kqh0Xvay/Qgyd1fGyMDXZrTXxP+S290
KCn5/scfl2ocU65yMqHCWWrkOMX/1qJjkjRtURe5hV2JMmjc/0drBmncbV0DSqPzJj6oi+qLaHmY
OEAR2GIoVSlRgu91dP7rp/C1tu21leqM3rc6pzL/I2zmFHFyLlXib/sL+/Y4hkmHLGbtM4oYRtWh
3vs/9GQmyZA/lAO14G3cy0avfOXmAJJj89h90sFaTnFeUintrnFGqRobzTFk1NmupKilnsqI25vS
G4VS7/KI6h6vPyxEGqxICPD2veyCYAiNVEtIXE6khbhiwUXp01yrIsH2fg41dI5Z/bfKkGLsLImw
kA4vLzgJRGgK/U4Qg8DBqdlvYde4VS/HfTp7fTL9pPn31bHZhGKPmZSpZRgPQvdO+qoNfeMHYRCT
sIbDoQ7rE61OAT8LK8jUo446zT/uIQ9Hco1KFBIzR5QIvv3hN7GuVplk3S8Is9jk3YyBPqr+CZQH
523idBoz1+7TaW1lHhk72e2uALC7877UpXwzpPeHA9CoVIWZo7xddFNY3SOuOVsBNQ1TiszcC626
aeQRLc56dwQz83Xk0z42RfwLlROMaHefjbQnMPwncCjtOEC524Y7d1kyl+c4q9sRVeM6WzlBZ2Bp
49mwku7JRE0X+YPwfKxj6yVYmynK4hZWIe3gLZPYIJ0cC4XPFFjG311pYTtZOqeNGcEXvzusdUkc
EXZQCSlQ2tr73YdTMhE+PEMpCDUHsWmC/1MuJKDve3tgP4Dl7JS+GWzsEY4HJg+3a/EJUpD8a7Zk
a4QUPv/3yP7VxwKHhU70cHWuggq58/yLMzXMYopcg9oCxrnLjPF9kZzTWubTBn3zhtvI3weN7sRA
l5AIBU959kwwszlQPIWi4a6ur/9+5/sPaBB8SqEL2iP74NbWixGaDgvwtZKwXHcvHQnJ9KleT/Qt
mJqDFDeMMENgO8Bf25q2XobffE3gEArlTXG2ulsHfVE+f+ac9EgMEta+6tdoLEfg/HTct1un1W8J
P3JIm8902i/00+BzENQORrQZ+zqgR2TT5ek/kZo/txzYP2fl42QZmIz8Kv7yhWphuAXs2H0USnJ9
Wj/xkrRNy/6I8EkfG4t3RBwNnkwYTew+QHRXA0ojDNyaA+SEC1TVkO901eQ7f8QUTHC1jq9QtA+s
YE+VTWRUcsUL+PU5cBFLwmyrGkffJ5X/dX/WKvy826i5hLDHrMDl0f+xKk+FmHvB3DLkplTAPjaq
fzEjrrlrX8/v+5yLqzY4quJBF4YS3hQs5LfWCiuMEhIG2gXrvJZXRTxb7BeO21y5x/9WlzSFZrDG
G+z/PJMBhaW2SmO+s2C3HWgdVESCcVN0qkfkCndZPieqKz8rVQ2ZrBBIYE0bhTNcJoC+MmnvWWre
F5rsKWKpgzFy4O+mHTOroFq6QclUnd0a75qFl/XjqUnTohd5wqBjlldEKN43JLXXcRBM9epE2fNe
+GMP0eUnxGy2klmiiE+i3rQCNIW16pqnsCbF/0Hk6LswpL/h7EIlDuTX9jgiHsdgvmGNKqWvtM0u
jh36fbNVmQMfZTvEg4TCVDZSxlEvtdUvJUKlgowZ+k1wkP4CJq6p6QrKaQNjf3dn2RdQIi6UZkg3
etjMvQ+yHqX4dC7pjFdK91vnf+IEGszerbaE4s/as2J1sF4sMttkrIeqk6spIl9V8JPat7TMjajo
YFz7EWIc5ulQeQx2Vj0PnWeZm9hO5ehvcLJm6LnS0tGKMHYW+WNkKGBqHh02K1ZKf9Rys51FO1tw
QHVWsqjNd3nUWKQMv8UTcJQCrBORdVAnwSHYwpvlHEiom2z04lZweXORQ1RstLfaNK7223NPxQe5
bOc6SwvtpzPX4LqOwTZtokJZ8kMA0jd6ESBasGq73xB2t5fEW/+ztOLsZmbDv/Tb29vMhiG3Hbmi
/1ywCpJxQ8FSZaSmuJZ4T029wlpejiylxP1BER6tXeltl84ONvMmV7OkrKuHbs6IUgaqDQFFqTZX
9rlv6P0tEFUVXOTsA+Ixl0Ku/Xcn9ap6sw28k0+9/fvFUTfdgLlJj/3djV9XJLzJ5VOqqCRYM/pi
DVek43pIvuyg1z2JjusnDBw8pbfNMPyWas5ZDyVEepO3f+2xpsx1oo9PKWpzjjwhTFV0QEkrOeEJ
yFHXhvqopZRzyC6IUe7azDhe4627OG05yEw1uRzm6JwXbfRFuaGbKUPmWr8Tr54zkfiuXcYp5WiD
hE4FaYfXGvUCLz4q0RhrDDqnklM1qAisnENtaMF0WfRDtViVtBFTo2a6sfcQEpFUyWXQuwDutLeQ
06utHLG7khQjRcqKZ/Xxe/ouCAcpyc/iSHufAPAG8Kcialg7kyBhsPThdHdIWP2uILVQ6ZoWNh+L
Ex4dHq+gWma6z1Vg4LwRt1Z/IaN/CDMc8FEFpK+amySbl+w6NI9uNTPlhTuTix1uihzTGPqnCQG8
2FHnfcxgyoIFbhX8VDLVcl8SfjBzLVJYcHNffl73rlQosN6b1uTRLG7WFWrCN509t/Td/vHEnHkO
Vwq/qaPbRBVL1BAY/+sCOmQDiIrXhSV/f8gkhuGPaXEfb/TRa2ObPpSsyG6Ol5M3XpwBh9gBKfB0
nsUOOjTZCuryUWzcU/F/iCPDLcsnJQXhod8aufickJ8vCZ31EWhKXHgLh+BTivFjSychygB5ZPyK
pOcEP560T1XWbJnIJTf4GHsVLtcg3oWmmxu81k/TMCV2prTJEaIkb+a1izgTU9pTbl3VVT76q7/+
kEKkPEsVpakcoKsomY4EGg7gFs/XcXOhwqSjntW6WWEyHFHv5HBttl1FaPSQwnWjmMhT0Y20aloM
JWCKZoACwulqPZ+FqN7UwHatWOrvcqT6uh0yXIXHPHcMITfa9XWeklJo/8VkU4kvdMpsouWcbqwx
+pYAUF8lgYfHVbttRXXxny0sf9OTJeVsqECjeMa2ShWoWS6HXQ7AVTDWI8pIm+V9fJUmiHgy4hbb
HhetFN9W6Deuc+1qiPacEmliVzcBiJGwFS9zqiUAN8YNGe29Olhjh6TjluopJpkX0Hgs7SFyOmgf
6LJP5Hn3f0JVQ5XH0EOJ5ZHMTHIEti+zJk8OTGHxdZAGDDlKAZTanbslsc4P4X+aJoAX34USG3nk
BNHfr6jdw6Ya+OF/+YkChGECMbjWETypZ6/oKrh42oM+6o9cSzzOKFQltsjZHqK01BY396i5OhCa
utoyPZYRaxdzpB5Kcgls0qDoAzbufjlU977c4STGKND0mo+1LC4FpGHJMpSS1eDNvAXYVGK89JU+
TYlv3F7ZoZTgwuR8VGD8cn5EC4RLX2yfOuWN0cwYJA4ATUxlfTsnYZZ2CT6Sn6Q+7kt+KQABGWs7
mPl26zT6lS8jON+uNG7SjcyC1HTb/ATNfIsSJfT4fvQ09f4SUdW9/aW3iZ5Fva32jgo/NC+5weA1
nDcCqm9JfN+VdOuZzCfDxlKGm92cFbTvy6g8BebHoi8j1IfSZ3byaAapxp6Aww+NPWDpL0agXl0r
x/Lb/RAo3YUmYxoR8Ey9lwc9IpiRV/QsR39qFCzeugwlpXJpW97RF0bZ6VYMOkoXMdAH9BuhUDLT
sk2EDj21VAY9jvSKjdhJEpLzBDG6m4324wXjpJIEA8jQ3zY+IEdohtIVOx1P/XbroAsJYSdXBdQM
0r+lvnrfjq5zHI5IC6iJJ9WRpJ0XnYyaqW98/+RiGIZpcLrBBcvJz2KCFCV9gVyQtDeMNPhPWnLR
ujUHKLF9w7O5/AFp0hLIAWCB4Rv9xvg0nremokHwv7MLNTA4M6kUB8DhwjNuNvr/W6kfMqLLSE2A
XeR0IywNBYf95Zj11tAh+xF+TtZ3lEcUx7msn3s4xz3vGYTcdKSFZ0JwJ4WTQym1RR2SpjrvhteP
0gK/nG/oS3ubPJfW3L4dzZzKNKaNEqvEjZ+YSz8U9XDtEzpyTj1aO8QaqLiBiRoENgocPwKjw+iq
/qeXKAiLI8rUBnQnTLVGkUdU9s6P5J1zpzNNiJi6xinisuyCcZE9aJ70xBMgZ+O6LWnf1/Ktte/P
hqU1/1hFuuEmDJy6VgjHIyn/z/7sofrQ31tn0q17+m7Y1PnuJjp3Ck8FFD2SIN7SoAqNMMqlHxQb
2ZabEmz5rmdkWnr0JJXmfHFYA4VJF4Vx1VoU8RbCfM77ou/Zhm8uER5sDv7SBdSQo4FfYQeHWMct
mQSyZoDtKpWlhAmjM6ajhnzmjMv5i4L902whE41p6xwn3QCFT5Gzlm++LONaZxk8GZgbhB0TrDMm
+hWWHb9wN4MB3i/D9Hz9QPxBk1lZF2ub+oguqvS5RLmpomM7yrVwrrhl4jvPsL8B2bRRqT0dLVT3
7jHXhM1bWpZE4Na4h39U6hbBB2wquNFK4U93OJQF1ur4YXudF9j4B70+m72GXoWDVos7qgwGrvkU
kp3Wr+J9YR0+WeFlfCPMplLvALOTS7qbXG5JepB38lMFgZucOnDbM88aRMHAY8bLvpQofV4YgDu/
5vFcad4YKfNX0xbbQ61gYTKaUg6MK3uJTLTFKO4Amw55/VcuyzaoQpCLqR5SHSjsLPlOjMf0aO/c
PQ5ChwYz5aJF2iV4MTc/ucoryP9JrUWF+mAphakdomDPx0uxGOduYLtdukCJBjA8PR8tu9UuG/J0
aHAvIdfof2NKAaVqlo9VGbC5qYe2psZDlo4iW43K9iEmZoHSM4rfwxipcss20FuF9IIdqBgATPXk
XCh0pTRB4Ttvz9GMdb4eevEELwVsKHK74IykgFXTNi7mq/fD6EJAO/q6T1HR+dKBxHsn13yoHSwO
ifzI08GRsku/HgEabNIAwpH6lwTVSGC7VyM4ivj3s3K0APR3YNKLowhek+3W1c3qeAINSCEXsQzO
G3JYl2NB4cANicSPUAbBcGm7mIcFaWvj3H55gRg0fLLw4xRHjn+YoqYA+uIcRw7fcQ9sqRASKmnz
mb+I/5qaKz/NoDVKR6Rm1x3TyoiHq/JDCcNZ0fhUDo7D3wl1OOwdZRqdmH9r2+CpD/K8AOVk4uL3
oAKJ3DeLupJQ47FsJ//JGfrbYuau+RU7fRMyNos4U0YMjw66f83cQSTtiDTOmhWs1IkCcHgrWibD
73i923hA4u0AY1WrqHglGJgGW4+4+R6Sas6xlzJtCOBOKgAsmUcl+LbbZK3ZKF0J7rWaFjgdhxh/
8F5/iqqqZQK3eo7/3Y1kpnDP7EWTvxRtD/G3ljVStS2bK0ckeA3GgrbWYCESEqE9wJYiE/kZpi7q
19faHExl5S/KnwgHIlfew8odvW6pB2aEI2/89XtaKSTRyNdxO27mF1n5fw+RwGb4hB4z8d2ykPxp
myRXzq62j65epcrEPU0qHyCMDj/DkGUxnSWE2xEVlHosjVSIcxpj8+0fwRw8QjMBKxVfuXdX8WFB
j46aoBSdQb+bL8TmfXSFcinzwWkEiAyYXtI8NZCDyS6c1gS3In3Jk0phJpmgVkyHDdgPUATc4Hhx
3jGPsTapYYx170ximvEixyhetNyIumHEjifniyeRXBbhrTla6x/MsqcXDNdDZ0PTrjW7+dAVAwco
LobqJrneC/97awPSgRxqQSNWAEzxdMlSBXePDGffooAbm7XpNEHbW89WB3L5t+9I8V/K7jB7DYFB
8g6TIom0jjbur1EmR/mq5RK9j6rfnUxjMDwUleeQ4fgWtR3LwYEVEe82nLEwktyOGjzw85vYWjt9
GqDo9ttlvz+yZmQNcd1q4vpL6lz+tnXKzsRcXwilYVWQlW9gKdmAu3kBv91Uh8JZzAOqEdJZsYew
c4p4UWQZkXlQ5PllRw/WaMgOyZ5/3JS42x82BsGmTMnD5QgkSDJ6UUJ6acStdLBO1UykZNGBxJPf
/rvcbE2EMZ0BM+Wq5OtLB0g/H3Qsg5IUHw+o2KbzKCw2YpQlGlo6WomBGYI80qpDiMCf3ex6w/+6
gQ7PDfDpls47qITfTzCcqWxB6xxFV5di4Ac2inwzTueroOWQM93srnRWAyejSZhoP6wS4qacj7B+
XCqY9eZl6t8j5OC/u93cdz9pEYHFnXcX9ewgvJJi2PJq1QRhWAawnbg7/5Gc9rQnRgFh6yfJoplF
GpHEpoxXAzygkUligORJf8IbaJATxcuXadN4FJdG3E9F6syWKZ1ofctzt5wz+BQfzavE5+kx35Lg
R0XVIwu1vlMOubkWe+RN/sMRlJ+mipFpoKIr0Uyq2p8GBzeCfAuHtM9lIorVsLJWjBVkqJRuQBBZ
DwdpYLqEVHqaAemxqAvwqojE0gDBNofYnNLzM8pdaWoNgTlEE2NasHJSRbDuRfadfi6ibmjiYDLg
dLMjY7HZuX/XvKV7VpajoNakbKp2C/zVPy49ihrlvvL7BLBr0d0+uo9H2hzQc0WiUvdZDSpzyL95
fZyRVgBISlu/UvECpcsYsxc7iH14AKqi11guPl1y5/Q5LYSWVMvIO4I0J41RGbO9Cszm4M5NtRfM
FbXi3VswUzK1Sa8kXF5Tx1qR8mL7NPTlNXY4LRJVAU3HtKNKE5mUPiIOpHxQEb4jDrzBBAoPZ8f6
XO923uRs0iaySBn47bGLmJWth0kIRT45KeZTFAjKktnHsXA3++jSRxnF5NJn5d8uqefvQJuA8gMf
nZ0X1fPefMA3ycBcaZSB9ryUMeeFSAGW9hy86q6g3uwi2MaKxjgzc8DQb/Mu0SHjUSF9ePHBgTw8
AHfLYFdD2m3BWsK78C1QevYg45+yrXf33tw7xxU1KeGsm5+jEDEVchFFyKv9IWryxsiy/JviLEaV
Hk+ZMjeUy3Z/5XjeM8jiW2B+GABA1pUUj1pQi1FxCwrwc+G/7xaJCYIHLcO835bJgpyqGO9j1qRf
l0onETXJR2946UpAe0IWKj6WXewbaiZBsGm6Po2HJGAc3q7t7PYw3/M1HLCnc06//Bs6ZTZ/rkqk
LcxfH5TN46q9bojjW1OLdSGjwtlL/qnaDtEVQOLHVdhMAIF3mXFM2/QAt4GgIXk0SOzeHElp3Nf8
LWavl3cJbnrt8ywICFCL42LWl2CsTp0ivWVrQ3MTn0Su5h3YAPpa+o1r6DaF1Jil+dUvGaBi1kyl
/e7GrOfx0zAExSlCXkKkj1jjxppZMS0ML09vxDw8/007mL3JrGKsmknu5zHDvbL4TjBDr7zznems
nLB1ZR47O6AzkTUfCDSEGLlLXzfyY3kwq1Mdq3FowZso/HTOwcmQzkkQ4i1xi9CThZCXu0LtMm7o
JKzRwguTS8atefOvFl9U4jHHdx5OEPMIYcCJJTr/M9sbnNEz1xdVHo62eYiusQ7J1YwpXs8dvb6J
89HAd8eBt9EVRNY8v/BnruyMqdoRzJUTeUCHZjoStzDAYuIRrHkvZ9/yLng5CBD8u1Ni+kmxV4wh
XNZVJoyyjPKMPQBMa8GRE4mAZdg/zWG3EbHvY+G9MMnrKKerb3f4VSNyftjbOjbr/9wtid83aGWE
kOcUQumO3ysWXet5ex3k8XLPc4dFdEXoLyBivy+ZIBLqHkAkctZQMEq361N1LBgox7wNePRxQM5/
54RYvM+RMvwg6rXHdtyGCr2MVbK+Wil1+62+9BZCKXi9Y3PDFn6PamcNGwzjHt2J2DejCeXcHMgq
GBPljLwbMjBb6vbi2IBDjUmDHPrWEbNHI9P+uiP6GnMUAR2Hp4mkTyctrdCqyEJmYEZD4gW1hOp/
UT7YImvYaJpsc582LIiH7nsey7ZU8AFRrTZoFq5ePyYBI82+Bdb7CrcTqfKTY/WkzGwOMexR++jv
3YhFb0A1BWnOp0M31fsbkP+GjsJ8PInFJr3pb8iplLORFh+m8SBv+lT6NTmnpfDlGQSUdGbg6ezb
kngUIb7lL9WfWhbv/iS/L2PnpQc3P4czfx/tkfL5Lgku/eM5FDRi1ykVTtsV1UtlPTAym6S4NoXF
tWrvmRW/tZ6RQCYFbkAFoKor6j+q6a6ws8NCiM3VXW4lvMOBsbnY5qSkaFB/PKYJqHbEAu1ULhg8
qrMIo0ClSMhrfMybTVdbGYOF2tqHg+dktmgzvixRzZNP5t8aFTVjKnW7fc4Tq8mRFbBwznkFPLP9
whM/alnCZHgQJEz/MJ21zH2xQODA1gKjkSkM99LQ2aykQGDJEtn+8O1kOjaVjlr4W4uijo5adtmC
ZlosdWVtVL645MvaBcwFGvfofep2HLJTOFJNGZ+XbgsSPN2St5THsPYJ3LnrpDfJ6UDrFs7WZzqn
5fIUucxbf7gsFqmMVri/xcT6EOKlufkXjjxN5igjqal5J3dvQyzit1AzPOu7310CPB8G/LwD5kz3
b/WqXGtVQ9y1/Z/99pkjUmvVEVIb1y2R43NwZacJNUAtYzwtj0pQuDzYXpgmkj4qeN7wT0NORvWR
ECQA2RBNXFA65Pvo7mfAPS1E6u156/R4EupYR4oIZE1YdehOKyQNImRadw7J55D8rcH1Xo9+IpSM
rqTxM0RZ8cqrdtxIllzGMzerWTcCoavzRFtR4MWE2vzEn9/dnsuL0bX2d+96qeqJk5QONZ9lOo1y
GdgGsh4sRxwVc+DqtKKGAX5+Chd+YzPBoihqLbLMObGpsScE3KZ5rhegx2puzveOw8rKwWPoRK8J
xxsxJb5gvbssmxhyiT02gGVRClUv9owAkxUiTt3xJSDcOs5R+5iinSSH81N2Se7FptEVTrPqHZd0
m9NtkeWW/4Ia49mun/kZK81kzN1I3uDzzw7L1o2J3E2hY5EKEmxUmWGJDkI/z+0XthpBrDT/ahDp
LZK5xvmRpsULP6CzuuJdFSNgvM8VUil8RVllMoms0vU11sz8KZhHcEAmdidqaWajHiyeEsAUs1SI
et4NefdGxd3P0VbB8ntDlp4WZZ49SxqMPzB2lsaSYLf9PH3zfBzEdjqQncPviUStHu9LenqPkxj8
Gu300W31MWLgqqCtjruIdhlGNGXTSn3vPYEf7QQMnaKD5i7Gd6A/nVy2WrzEpnZh1a9lb4A68Ljm
YQttjKn2sRzsrw/isKEHbwIBXdc+tR1vYcDXT4FC0apgZRQLAss3Tbb6L3Dy24bIOyxIac3sQJb7
4/AZGG3IrWE5jZAU1WQ+9XPqAiiwMdv8AZfmG4G3HUPykpKcq0ARxaLGZPVmukRNR/zh7KbXEb2w
G3XmqntCYAeyAp5fFUeB5lsgJQfvoVeTaoSTM7mM/BWrxOZfcTvl4HZWj/+YL9jPBxd3CyMJW1dV
bXtXPnruovKNSUzivygXxcJ0DgSe81es9Hzk3ML8hahAGKGZViQXZYF7px7lNrGQNSD6hf6cw7bu
OQWpS46h4ViKizhGPbpnKckZtFxmZHClpvTPp3JgWHXLhOINO8M4Kc0XbANhDUU6aqGJEDgEr7bC
EbtHxsMSLzmjHNkNIFI1vjukUt/3F6b8i/dVtdV+ICG3RJJxnEB6wN+XCLN8Bjh39DKVcz2hU8As
+0Q9Wl1vIIoPtLNTfQvjHmuNfTsHRTH7AOvJTDzenLJNS2V55ICc4DZ3OoZy4vucP0ap7iO1qB2V
TZE5AIACyNzrKo4BR0ipveqjO15NqPnXlomoxjUnnC4O0tyFuCb2uV2sQFaq/GMXK1mAjeDUaY4D
nF2uTj6i4QwPqfH02f5X7PODpSHltQJc4FkF8WLojNpS92MTOVleJmB5CL6t7uT69Bsk1oa+X1EJ
L5Eif8ZSvOmoB7IgAIdAaRJi50VgCtbEvvsaVOO1owY25PEjIK3OUEHZ+tkpANapxUVUVCZWTRB2
yd/qtlGzgJA7jDhJUqsyupoqO4A1+QSoUjRFVQ/fHqUUtI7ANiz9fD1uoWbRhEv1NUa0SpqkCcvZ
n73EGsyNXYTOeSJuzjWuraJ4CX6/d/EeiJaJ1LJ0c2kd4GHte6GCde6dCtbo6tlgq+od5fNWzuE9
1vD8D0zk2HsksBgCWbSWH3rXUbOsKgovh5GEqKYue2SBEuX32UCRBn/uubiVHiIb8XYU5oN3eoGR
L67PWoGIZ4bkQ++zjVBYqJjJy5UO51ttTw6y6qolPgcr7vetTvWGBcIQTFTTVE1b/mMqDavx5+Qs
RqovPeavdjn0SGiEMIO7GK8ovWaTVHbp5Exnsc/CtkpJ1jwVlLMxw5fdP1gfxXf4oX85xEyiHrNo
ueHKXLFrYd/20mk49Xuu1e2qbP1cLfzZA+mf0wreHNFnEYxgOL9DMrsbqUv6D/DSopoM2vhifNfZ
US3mVTJGUS03DqPI5RjEACCew7Is6IXzQEVRzjVPd/9tJFkzylogQmGEM8EAM8b6cl7cqlHEEJa3
wj5jgHW+ttD806UzF5UlH5vXW7MUwMsUkU8rzATN/SOvmmkJFMQDSicMx51RiyMyEcjz4e2F/fY5
S0hqoooFmOuzfhwZgHgzKCm2UG5x3KWiYA+bT/SqeuryYaGqQhTTAHrzRjpbRei+bOPc4Q5FaH0L
5cIdIf9qjTv0JhZLfQBC1HSUffBtCLCTNkGKvqShpyk1Iq6YngEINrpAW35RlIRYCU39qxjzb6tS
63f9Fi/hBVZyGR4ziTA/OlER9b0npiwNbTN4fu7A7ORD1DMGE37I62my2Yue4/Bbqm+6lAQ0iv71
W0SEbboojBMnOdQArq1JEOWoAp7AnjKlCtr/XWxRFvTJfTfQdhXR5relFaPYw4xjavxOlxC8U+X2
p1MDYyoE1rb5O4+G+2eXNvqIIGhc6GWY5vBqM5Uurlqc+9CMDmbUsZwHB1gufo1Ueoabw8PVxjiZ
l5xUNW07qkZDitIsMzGyp1eUrhFlKVkLFWTSRdW0pHgof1eCe6yYKp+Ypf/QGfRwpTeDO2dkLl/C
MAVqNXXXGA7hWUFoAO7FXPwD4bpjcxA/ijAMVbibmyfKe9okXPbCRIaQ03IrASkYkUomylBJUNbf
f7oZD8yGQwdd5zrOOTtG8EC4hTztrdVmymr/IX6zwkRUvS86ZG847P7H//3VepKeW+iR2m60TBVe
JmJQpEzGi4/AUxg40hhF7qwehru93EjLVomk4eLd+4aqX5gXSriXD3qGicfJFGXbeibxfhhBzh06
F12XL7Ehts2EI0ze6pgHsUtX0knHmNSp4QKNWHT0paLYNzmTI4uk2UEMJpXEUamRPapNAMEpOsCP
poJSkSfjXjYVIxKBZyYzjSPzpjxdmVSY6ycm82e+0Ekk+ju3IEpiGeN88oqu6xfncSkfJmR9k2Qg
vT72y32XCXhFGApgiNKh2Bp8r8MXfr/nWFFTtFyJ4K4dhsI7ipVLKbIUSDNbmigzaa95PBnUVPtp
XakzTbzJXr1JCxqml4VRFNrPE5i7NYVWjBfESunUmEW0UFG+iigLy1GZ79PykyoyTs3NN8CaCm9y
lMkOii+dnX5OsKM1bN0Gq1HWIigMRoVgHFzdZ+ZidCQqyvAwnNX5mf6O2VwVwlyB4dPZXjhKDgzy
mQfxfLCIFftJw3OucC3zSm+4VybPE/g8y2gO8DGug+0IB6P/RKAD0Ms4kxD5ijEzYSzmgORBxrrM
eesJyRLLtDd3/qzL+dvXYJpn+YXp5afhiA5X5q18WAOZhfQm6DcaUnISzWUW3M/JzdBK1OQxAvfO
UBXiyjOZOSPmhH+8ApwSCUw/ryY0vDlu8WGQurXpbeiyZZIDGiGOQ50hCv3aPGlGwvxULkXsgRat
s+WsL6m+ZLV5I0IaUDytc5hm4LOZXrZjy4oPmLNQEStUNMdq04BDnslmKWuVdivZzy9icEupbexG
1IOozdQ0q8vyKwCKrkUSwX3Vs5V35vyKwKuoEdDhwy7EWURgVEPrpo2/fprtKidH6bf4NSWmXwZd
G5tPv8fk3B9dLqPbGJrsQx8eb5YxFp/zNg0JSXQcWCnrZ4nYynMswCa3i8yT/38yvSAizMX09loL
tFzv4ocRT80vKhc1WqoWFi2WThpT87RC0GZk55U6BDsb5wf28GgRGQ3qtwfzL2l6gfSui4HY/BCe
YDIlV+f1velD7HW+RePIa4tCqlTjIeJn846fcT5uSRC8lQfA4pLPDEYquhJQLdfIiMphtCt+hDy8
6Y+emDe3SP2FkrcaFh14AnSJg1H843/b9GkIjQJRRMWfOR+HoJll/402rpJdhYPF7jUuQsZZJJmO
c9gVLg5bYrh0Lqi4/1aduFEWV6RDGULwxJjyP9pYU7ngzKFz46QM5UVKi1KcqLw9npLXJVINkyLq
1wxmixjCvRniv2Shja0shLYEgiCQp6EadOmMkfSVXW+33QiTK5d11H60a0hyZovYjYd5/Z2NlQM/
olnW2e4sqYujd+VYDcv34/OBG2q/udCH6aAqsw8MvML8UIlSB+FPxEuWE6mOPty4zuLTTNIhQxEk
PuGLeI3YrSRWgu2C1kuWKtsfghgRp6CUCRyOIU9qJWYHnjMH8KI2YZ90lMEymq18qyN8xuk3s9SE
WWm8dX4C2tIR1LrUNqfhSXahSjDtDuOpRUKfgdGHZjko0K/Tc7mkLPROWyDU1wKiJhyDpGSRf3+O
3bc9PhSxyAFSlqiAziU/xf8mE+rL6YIr2o9hmb9RCOQ5/AED2VcrCpOtbhVU2n50HgStoA/4/Ask
l9N5cNjVHkc7jrhYdGLr+aYkkI+XETXd9iCtEgukAgxJ0RXbjm8+RjO6aBHzBqOUehI9udV4Fg8b
Ec/9xguxFDtiWhX1WSwAjT7qrpMfExepyATFJQT/sieSAz8NUgSbE69kbGGaUvEzs3My2j717YAd
PeYJYedfeu7EM8Rjt+9p9Cs2DypbTA0SyYyS7INsyTMf8XZu7JgtJOHh5v9o4fcie2oUOWc4IV1C
Thz8di7DsO7O70FodMoEazxr6JOVa2p0svsmPmLJOtTw32C4J8FbxHecLx0GB/TRZ6oL0tZQkcNh
Sd0EpNAXXsBXBu0ulwpH0XZDxHzGXB7GJkj6TMXj4wrtL9eJNbsSRYFevvDTe6siHQ2zErQR96h1
MqJot0Rmdc1vmLJT+rxxlcqdhp2zPc3H9ckSXOxd/98IsAktuD3lAiT/j7oN9Ctt3ugzS0ftWqFc
VPLDMMLC3ADBWUskXYjx7His76aLdc8u6ovXORdqNLEypObZDEQkxuwXwji9JlSR5FYhrQF9blga
kAMnN3XjBcyEPq9A50FThaceIsPn5Ve6hvHVrc16uXHj/ROMWSh9s+xIPKO0gJGSXEgPXFCby+ag
BMlMbqUp9EkMWAmtfXK9i/F57G11wUbkE1+adRSycqH1lkb44vPHNRcSE5eqHLIIq18dhrsQRnl1
Y0dHXjByvOFPdUuzB2j1wUwZD73sQClan1jggH1AsNzvAmr3tjNVp8dmSRwGfSFP5IeOC2Jfv25W
bcNMsgUPFY/sQQ1lC/yJxnFYLvxUVZY4mV7xeuwvhdAFqCItOOwFS2FPAtuUy3KTjkm3BTrK/xVv
oUAMsm4lf8CqWJTXfKOymWNeCLbhXyafW+04bUbbZaaAlXfIA2V9OcBA0rbdlgH4UVIcI6LPB4dZ
GtrbkwOE2aP7xxmVYDxJOGDEuXFV1IXQ8kBFa0ExK69h8UDluk8TVhiC+OZNJLVW0JXCl7pqbUij
TVOeW7xcTNvIgyOLR469CtJxdsCsgrOAzAaW9/OOt4zUQaRHhacrEtzAPznY5syO0J1/+Wa+1LhF
ir8g05P6wZ6RwGzgBerQe1Gxy20QPDXvBYhdHvAR2o6LrCntJK6uhHOuFnGSmY1NflYoe3j5/UY1
uBDpWFixCJM8RUAYh6zoiWUkgx0wwOQuB70aPgWcbN+0tMY/mCpIHbQoLXCtus1omTt3a8dFdnBt
L/AITslGfJmt7Azd69OJdAWgQh9mIuCVGxzoMO6iYlNHVuDn7rXnyEEHdPLtYbJG8tphu5heMkKJ
uaiA9LIfs60oNrpSYW0ZAh2GUTc8EGWbtf+sC3m5RlApZFjQEsza18oCxfBPf8CTlnfbDWVRKYG0
hmdAM5Ut8Z61zqv+lGEyb1s+TnQNLXLirG0h70eFKOmiL0guEzzwerc/DxRf9RWU/b5bagP9VMGu
D4jLkJLCIQiPMYE59CjiW4QL705v4734gBWYB+JCU/yYLXpd7Cj4IFJ7GaXW41FluGgLnlFaXDPI
u/+pTxl6nmsIsosZ9UMpSK58231q9BLcuEb9wWLKr5pasPLiquj2d8M4DxlF+CMD0R3PXgzCqmvT
Pyq/f7pTFHNHTcExVC/cTYYsHwy+/bm08nFt+rP9D6BkgNc+qf2d2yOPAsvD9IEwCS+f1xzZXLOP
nend8M1YXU9ku7b4jqKGwYe88EhnFSTjwt+s3UjHY52lflu8518ZsT/Mzx/lZQRTpyLRo0+tzFo8
F2mB6GY55jPyW9ZMpL9HsOqtffRmO7DWBuJZuvk1lBSeocEcFgYDKo8RCRxAk6YZIlOEUTp0rY3B
wBVVxnOgDVl5/toYYdink2Tsd3wclxs2aWJ9vtdkESS8sdXw7UTAwWIVZxc6jP7r5+iJnzZvzLER
UMo8HAfzsPqGwEXiymfuyNYLhPXigv2qLcMd9s5wc7ZrSG6m8H1Wv8SyDbZTdyIUSBpJOeo1rPQQ
61iHZFfqg5UM27JyryOn7pEM4NVpTTEkQA0hXZd1fkFhrtV9xtj2nvKL0j890R0JLTz3Gws8WHAe
wIuQzCdsXLpJj8J2igbeen1g9PXA8ChQYT20PdBleu+B8E3FuQzzHc18ZV4r4I0T3A3P1NrZRHQE
MmSMP+xnohmBd7iwgpYirFel7FPjOKKqNMQ4GEyYD3aVIcOFlI0JYe3mZKG/ID6xnBA6y0g6zDf3
/UqPlcYWb0MmsFvfJIEciQE1ZZK6whZ9wvftMvKZLScD+B/nWDszLUHvyZlaKKBCgPCEKv8Z3lXX
J08+An/C6jLg3Jt18BY7IEp0CASDdr/Cyuw1lEwT6YOonBOJnNNvngkJXQaScKVs+4zAXy7qu4Z3
t0haVNwIYeXTjH+IiK/lClg66zYC17+D0KAofNP7O2SneXlBaI2csKrymv4anf1UeVP2QI9u4kPw
hLqPK5DXy1mjL43OX895qb+3t8q+cuJKs2T8maf+Fc+NYALtkDovNFEo/J3iPZmtRW0ePFjoMYi1
Q2nww18Uv0dxBj1AiH+ZIIAJE9GfzPdE7tzi46LldeV3V/uHJVDJS8heIM4PXWyZ21LiMev1zL5o
PM04eLEb+2cjbTvmKwLjDN72BkTFvgJ1MRTfLCL4KIr+ZCzexqAvkoNjBtaA2Kk19K1a1lbSbeGK
OuhoVRGkX6fPJZEVt7LlLV3FsdvFQK0+LbkMCU60Ccy2QdhOpS7MiilGRSyHYXeeNEDm4mlF+FWD
Zc2S7oPhssauQc3XSv/8rl8s2dUEHAP7M5QDUtl/AYN6/ZtM5Y5AQjdC478kTp0fPMJnMZ2sa9Ne
XAczZ+d+Pu7LUjqjE9IT5rPNMrHM4ab3K8JCGUZ/+a2uzpA3S6s0Vkl02GVxtPg5SlDnYh93CFeX
8t6mrOSwlHJ2vhuPymlnRrqf30NCiTZt6pJtIx+mlmGWsVweV4qB1FXYU4E7qzjTY94py6m2Kga5
mCrR2dKOqFTMdihr2Rl4ptA3iwGDQchpyYI70zY4Jdjl8hm5OO66QaiOeSgrHyB5BepXklXzqET6
F6TE1TKz3t/JnpEnKQs+iGRVrcprVIvLvUQ5ap1LeKqHVrANmytTy2QBZMGJ1lCw/g1Auuu5LXZa
XYqO+d+2Sv1RvoVbLYBARhTTVXXiW2a6ram3VIGFj+wVg+KI7EjxvxhuAr+rd802foyBzQBkZsfw
xhdVm3ZBVSuQ7pEjOSVNcUeidS28JO3q5ANaSqJBlOoSHGdX4sflLVeaHFK5zHWoap14kFGReFwm
ucbo9KIFr6eZXc/rWqepIiQI/bo4FfDgETtEwvwyBXxyHtj/9uuLaosoK+/XM6n6XnUXUDDo1lGf
F7qzaVUdhdUJNl9rUhlbQeXKeeCuORAdxQPEkXajbVMpimd/N39ffBwZHoBnQ6PAODq4IRDQ5V7x
ZppWg6lNUvlsm1xG2EFT5PCwjT2DCr4Q4r/5uG2vAjtuHLbpvoX6bExy2V5daces5sE8T7vzd0GH
+JNN0PvvH4Mt2UD//lIZyuFPKGibSo2iSrqeen6gErE/tBgC5/0BExAsE88NkqyWdFfZa4RJOFv+
bxT2vDQnOQQptQFfe+QjfTKZZUnsKtBao24tkoXYgHgDOJQcAgCAoGXRZ6/fAzn/WjQuz0Qop5tc
EpOZWCgmJjRrAYv0VExc/vcD6/opA1qHWvJ1vfRTJPnEkxANJxBMfMNgofKmiOCmuIDNiqM/G91Z
K2flDcuDtgG4OTapJmjmlRuQSNVDxNCfZe5wEFXOWB63+cahba/xavk7DVHktPxgt1A3tPkA4C4F
M4R4/vjt8wrkfWc6BjlM47EP31dusesGhEsPlgnmlGDePqlo9tt1vba/LnZhhI24BOwhrBOXbwRR
0yXpUKfaKc0AfXCGALJ3sltUCvDIcv73LaNQvfVlGpaEZUaYd2b8ukQWRBUTwdyh4+fyWjXbUtCg
24FjWEKGfm8vf13GgvwTm3j7WeWrNw5cjAP6ZkTc4G72q+C937+hOPEm58fpC+ivtdHgTnHz4skG
/YNI/zwnpQH72hAWIEqTN0L0AZab88iT9lPjjrxZLSra7NzdVAdgrz01fvU+e06KGtNOCd89pttE
kNtHr7Oi56DE7j/uD8xm5o86snS02IfgRCjkjRXFmE2cQHggHHgQU4FsHjzc4YBISkcMkQ4RWubV
XhA7ej1uhKVTq1pZjBmRhrSqD59Opgtfdmci6VQyAz7/B2z8HgLM8nIo141/LmlFHBXOF8I+/Zd+
TAKSXHSagRcTyQlt2Oz9YicOMP1SYOj7qcNrn7xJP8jE0hJVFqHYYlAMkNP/90VEnIRdo1ifLTxv
cI6mjiuJvoJrceQSW7SVdeF7Do7nRoGn8z+SxoL3WK8x61830KCXh9YgioAvNvavTImgzNN1BE82
oxf++gGkcRFK0iqcGhottHnddVC9KPyKeASYui1FArlqSYzkIGKg0izcT1NqVAc3NlKZceRs3j3v
PCrqnU0tDQB+MF6I3e/LWhC2z6kGMXKIM/oFCLt6ax8aB2sDquuV+jx3Q+b1dKlQHG0OdZ3pTIK/
A55Kprz6Pei1ujQ26757bmIN2PVPqy60l2sFZIOxL3KsNRyxHWJ/ltS04hTyGJa/FPy/Ljp4Q+Dk
Gsnmeq1JDCIFbYHPqG017W8gYtzEZFqjcvtjEERwQqaVoqqzXAQwKpoiYMGpvu5tWAL7UJIhoAph
EGjGJN6HeUMpGdXnZg8W3SD3Kx54OuUaB8M+2rJTsUrXO1NWrLHV0H5AMrmnBQEJu+jnR6uSSmdW
arIMuusdRtPDJe9OVMqgos4bHN3gDiZRMI/aVbsbU0zZhRNUYkI5d18Aof6WeeeNdQF2Kbfbb3HR
9c5l37JK7rJrmsKXG5gaf+vRuxo1Cd1QbLq02LDcP1DFuczrSUgmvV2zRyk7EXSkCdeXDU39/9zx
08icWZzgeSx7v1CTHOQwzVxIheuOV+xV8a3fTFVioUJofCGuei3lpKpMlmn4paqAYwnirBywGTAW
jQVns0nqQsfQtH2SMw6vU6MARSLihhE5o8BwmVtUyKhZuOS3Gtokq+dV/iTiXSwjCv9Gq53/wZxg
tk7VgXegbbb20toIwQuszER2xfH+IAgNv1qtNnbtgvB4N8u1k1Yu6XdiT9qH8qhWcjno9/rDekDh
OKX6MGfElcjOSI+7+xGBnXGbNP+ZeyflpPBUTO643qIFGRgj9jk81Q4alcfaENecAsy6zHvAD2dY
7mNAMRIA5vQPzscKkC+QbhlzB9qqGXa+Ljb/klBIoAc4diWcwJthlf2tEMASVWlZfZ5K8cpq0ETC
5uhy47PjXEaipwyq6vtHkVWHE+F5qhbti8RIpUWo3tw5BHTmxA11aD5EzzkuZcXgiYbgMpNKA9Cp
oQ3cnFeokMiURnfHrBggM+7/wikAa+sQlaSSi4WBIoqMKfu90WL+03cx2yPUQHlRma2mcLnAP0Dt
YQ/3aRVR0diEFd/JSwk/TiPNwKtcenYH1D2IB7+jvejRAbtGyOwacNnpNCdw6LQW1ul4gQB03v2z
bjd4VLbUy0sE3q6XlcWiqNb3GEbqqtL4YJ4RdaujlgK3iGHuqaWFeOQduGWtbb3V+On70hrCBBVg
pUNh9QdAOJv8qKn464jvnDAk58pI76VOtBIcQDXWrffSMKol5rm2PxIFbvbuGabRZvO9WnozBROw
PGAGXas+SBV3hvGxfFEHr6ZlB+s2T8Kk94L1RVd0GQoapmvLk3Mz1SZe+cnmlqUVT6eEJJatpYtD
N+EEBc/FQolrZLVzg1NyRdLF46eRUzJcmbJwMpb8rkIwHOyjLeaiefzv5Hg+u9PASBbgEbwhisym
jkFgsHUmpZjUail2YrXLAOk/wZBtffziex8wM8hFe/LvUpJth/QbCalxBPvHmOe46WmEBQcsXB8l
0HiXC4urKpawGljmkrWSLJ8pE3pNdTneaIPro2Tbcw5cYDjnMjnMFgHLOvnWOiWLgYCCP6GGfNyW
9v4GSKotSEs3y/7T4T+XOCyw+qQ2gqQDjmKY1gRH2CdXqn9TobiGZXb8cBRvvOze2spQgwV1HVY7
xdVP2smWILO7oFE81bFhirCd+gaAQgjQJlWYwuzpHEVAWRFv2QV4MEmtSbFUUhKGOQo8OzCYyb95
hmld0K8mYsd2MLmogScoFBMlNIPCr7jyLeTqS+KiVC/JOv+ij/kUOCgL0aq7EqjVkcm0fpPZDlOE
95YTmt9aaL7hGqF3fDZMOW9fVfcStSgeaJ5AfmuFIzsPuC3UacrsIuJU0Xcj4CL6MiCAIIfnXC4U
g4IaXxEyq5VOLKiIibhIB6BAVahrW6kOS2Jpux+6CAu47ll8XPLQbQBCOneXlLtUdCcWLAAckS/v
pxqs5dvtHAk+q0wsN0+1e0zeHjcfEtHaqs8gGCo1jsWG+q3XtLZ6dYbwJK72tTeAA532Tvz+oMLQ
lAaBBuVy81GOyu0ucS8FxtnwiZcEJOdog63n2WA9zMtDjKmehgFn85Onxsqx4f1k1mRW6uc2vyWG
H2wxwAcFf0ZkVhKmLPGmKdHaJO5alpwBsR9dfHGEm5eZ1x5HHmuYZg6wdYbX/ci9+65BHhd4VqBe
7YrskypVLqBZpov5sE1rahlMu4Tq02ert9p89XI/0EHGCuumGr3uBhkh/o1iMtI3xRtMxsghuIGE
S61YBEkQ0mNkC8s7dy8PdyqzgaOh8hisYt2wGTGkovpJ7qTHEKh28Ik5yPxLrYX296RIWskEeQDq
c/ihTuBuNXAzL06nxX6zRKYOCJeobjQOc7xeFvhdsdXSIBezaP1X1woSzhD9jspK+WzDdjMqpwTu
065LrNYJsFzOYnQj0XRL8DxLJfTHbnUexzKbu6FG3YMSZ7OiSWJ6x2yS5X541SXVPK2zDJr4iY2k
WqZcmZRgiVClph2cr3H1RK8YMMHu102TPPzLvQ8w4DK0UOUUZLmk202UmiaGz6IbRw2Cxh6mSlsC
oCnPlRTUWnlJggFbN2Pe07omItbHlU/jPQsrwuhaX8nu9094baQ5teI4CF+/xc/Qrq1mcfqjUlsj
efDfXhfJclT2k073OIwlUm/WN84URyqXNA4nh8Fg86+/Bfa8YwoC0gXxjHNZfGh6A01fXn5h5non
oAve5Qq3qyutzniUbVHpir+At8UbpOJiYr9fHBxJ/ZmJG6nXNw3a0O2jwdNK3JKypOBpoNRpVatP
vFD9+GJQdMrPZtEkEoWSBMFiSB3lgblO6okt9WB20cwzLMMHU7eQmrmxPCWzjNs5ho5/MSNAoPtQ
djvHXBVzd2TtteN74TfnoeeLGFz0JjUuo9pqwQRnkVBvw/MO4XZhkAdYDxIgjQK5fto7G4lZ0N/d
PIXp5xZSZ3DBqk4TdovPn6EZnpFSYG/Vg+0paLHpUh2XPiaYTFEUUhNjDWUEuH2igYXenWJZnPsa
z1K8VJ85ciSto6reg+dOCU0j0zEicev/fKESvl9jAVqNGhQQ3nfCgyuh5vfWOtMVWvhjtz3PpsS8
7/f0DLXhD7E/SzlGZqSluG+/relmpuMBkA4FT+qmjT3v9YGbpyhx+/4Tn9uuWxUSzb/Q20lqLqh4
zxPmo/cIpy9D5ZeQnOZ4N29Wi8GziKevNe6AWSRFXdSMeF1Jdots06GF6BAXot2Qmk6WLUtfZyJC
g5jH3AZjzClawT2sIV2Fwyv88Zh5bfQ4i5Mkwjcfn3sJoarQNuvLvZsPUspznTBhg2A6ZTZJK/v1
ihxvgmpAgCn6hgvAKmztkA0kORq+g844eV6ZC9nxIvr7u9AaIW+oi8mhuFpke52o93uYHJS5DaSc
1Pd+DCDM0r59JIyX0oSIdJtuTjLMJr28tbx8jyTmUm9iIX9a/wmpyz0VLQm8UBSPVsVJLFSRLxBL
re292ptj/KcTdK1wGYetda6WgxTzIL/vAdtFxJk1JPqyqt0vqYdm7yE4SH9N3mUvz8rMRLNPxBph
u1G5bOwfu4uBTdu4r7jq/9XJCTGVSKYd3V1O9fRMyNAOuy7z7h8zZUo6Lxna7sq1DWAbDqvfS9T/
Q2jHb+Z+tx5n1ZmSJx/elme/FWwKs8bp+XYs0WEtRlIN8sn5CEQT0EFASxMUOw8d5APTcYjTjjyj
DZ0XZqIfqmShpap/yALiVKEHOwqDvHZE+2o5owW8FiX4qcuuZWOb4Tce/aHm+aoVrmTQTBGOULUX
4bD0HuoZJLqRIZ2njJmEkpUPypE0mIIUIQ+g/UFFtlwPvPg4bN+fFoNR2eYoWpkVy25tAwEQR01j
T54D92UEfZwXr6sukGkXxbqzgOpBwbNPCLdFvMAJqITBFBHT7Tz5vCSXURL/cwNBT21KP4Aqz9nc
Uoj/bph6qpJc89nsQ9hqDlfH6+kkiJfoiL4119SGBJ8qqcTGFKkCQdRGiB2AUZZgFmmSfeZuippx
Pf4orbIyqKPSd4URCiiTiMLsfQYUvXExd7PumB5AsdF9uDK1dsUguppvscfwLBZlh0Zee0oFwiFd
HRa76x5R02V4F54LdfFzKZiOMIAsnspd6HT4kZAD+HgC+82snvkORPRxMkdicbM8ow8x2odwLK9i
CgJv02piUthOfUOKdm8JgqCHTV1WPkS+B1+YH7ps3OsIZLmGetsWIRmnEx7l2KrDokW3hnDZ8G24
IKV+angFESWxnlS/fARGRZEipcs64ogmYS9n53poL1SNr8il2AyRR/0dQ7AjDghdSYDCtw6oWU6A
6Fl3pK8UPv6wWxW80XQW8cnL6lklzm2d14HKpGUfjhWCCo1Pfhf/NSsxyzm7xNzW66vFn1dKxb2c
i29Qa5TJlOcdvlZkUW3yeugZvQYRR7Is72y2xYvxQzAKJKmyMQise8IqOQzhqguNjMJthwAzlRtX
pSkEAFQyKgLF4yIv44AatzgnyRDml3Ao1Wiwf83gE0yKDy4SRE34ke/OntGdjmGsxcIudRe0nQl2
yhmlqZHD8SK+QRP4rFX8kXmDlIYcKKc4pK6OTfCjPW9SlBFT7cWmIdNPkT4Q+InbrvE1aWDOnw+6
07c3wp3z/YIfJbAlr7Vd9i9DkMfi18tmHoWLBx44dNi++s11J25Lme/DxGWS8BCN6Rnw0a3RPUAc
FG9s9I+xfGR7TvEmT268Zw52iG9yZu855qge+wKCMTI4Kofn+SNCZaBGuOJw/ACLPgYVNs0YpB9r
ext6IweYOJJIm4Zqmf5wklBgVbRBtE7gUpAhG7rBL1WVQ3i+eaaSecvBe4NCdUWSMkfCL83dK0PK
mTG41+2JZeuhk6l/gUH9tXfeBWp7Irv/I+SImeBy+FRuOO+rnxGX8O1NphhkyW+rEeSTXM+KHcNR
zf0dl2npKAb/Oc77jUCsEcoBAyf/1psxzg74sBVNhg4WxKRKxKBTqY1LDdfopkEYK/eM9lUgprMi
r783ygg5RISRrQgJ8F6QZkWdc4iwQFX9EHlDkX3LjaNOkFBdNlTtxMY1gkpeZOw8qovO2moJWG6z
nvdUKJyd05aAvGvoM14jZULtK2x+fa5csvLovaYMRqBdyAVr8ZMxldN05yuNyDm5Yr8dviUEeC41
PPPYYikoOkciEkYazJW7vbPdH3yIzE9THJVMZGpZBCy6lBNWmj7NuEtirjMNqyriFqOvn/lKwHod
vceQoaNFPhFe/Ikuca14bESnw5/TVqOjdgvMAzKWJOdVXHarZ/TZA3iWpQsUskJ4G1pZHKDLcQI1
fCYpGwLJgxug9uSglqzO6oC2o//kvIUwBKpUZIqoJncTchL0Zb4r/EAgIwt7yARpTbZPVOPNAEFi
gBDsXxwkgkPV71ANRld/K8YDGEulHhdC6kVn76jMoAStjSfs4qshiEwXo8ARLWBoPlyBkSC2ySFD
8lPeFNoFHgs75g0xYITKt8ZPMOhhMW8aoSmVSmVqmAdDgn56iaT6t8u8XwW/L22WQUgWBlGv+PwM
p+bM2hEqv+DrVTDrPY/CLfvONiIYWBMRCG++SWKPZpRpraTvhNu4Y4q83FH08WByZ19lXBB8YsVT
h1WLhVzeXVNXz99efDQCipC3wQkPK4fxLI9NHDIdvFjZ7o/AU/19Adfg2P/w65KdZEkdwjRsLNJ+
5WHutusL9Rn56CkMiLrXiziDZNyzrgr0sPLtxpQZlCE0f2W9V6Bi/AoUMnWZyjNjHL9nyLrhPyxP
PrOIg4aBAo4A0gtFd17jfWrdYIizDe7qc4XnVDaN53LTP0WJf32VWcxshAytjD/Fs1z+T3WERFYP
ftiGYNfbTPaG+UII1M+tdWS1eVHMx+m0fwCnbwN6mZ8FPzUI3i7dXAibIf7wPbQIsoIX0zgBGsLm
2TELwQocIlbBe+OE9/rEMfRVc+WtWnbkJl98JZ5xlOV7cqZDCplSxNsbu7ab1QFUUAhaNvr5qumz
ZRi880kXJNxGEmjS+OkC6QJzOnsgKq+yVEb6Cf8BY0ZO0K/5+SAYEiMMr9Rqe7x5v2WyQdTuu0Xk
gK1r2qlcd1YkMm6QYNHypsonLEoUn09zsN5xk8yz+M2wtZBz0eIVGW9+UR3QQ+r2IooQxzal8wvB
qBN0ZOW38qNPHxK2gb0ByVEfCEVOg29IXnN/Q/7ziiL+6bIs/r9ojsASYvfRR7/clijnS3wfZy+N
wivJ70MB+jj6KSTEpy+zxXG92x2H0t4Upu6Rwhti9V3ws+48GwLA8HkpvRJg5uDIqtyCOet4c8bZ
qYlxGm/YI3iwF+hWooyq3e4MO7fVZllf49T/8hAh3lH4X+DVgvKyxWptPuWJ37K4zJTWYS2x1Kst
5x4iAA439h7YeuA5Z5ND3fxJ2WGLb+2K/N46IkuRTq2eLI3HXf8fOJ/p4h7KAxwk946ZrV+ZRSBO
JSLh9M5o+BcIPRbnkdG5X+B6rt6gt15adGahBjuC/rko8BSBtamAUx/MRjCKbRDY5W9GIAYY6ic1
SZK0SmCKXhrlWRUks/086r/R9u8y+Pt4TKI4BYjjKUUVgJe0Ey+6bN3T3ph8ODb+tHHMQfxfWwHN
ligCwmjkp5lxHm6Y+NjVCu96PMZFRLvh0HI714GOW3rYnNByLL1IaKtyR6CErjBisJ08tY0lYvSN
afgV6E5NvqjjwfoifMzlGi5LSeCFhgKg6Ys/qvRfrOTNYrKaSHQ0u/SgYDlYdidljz6fttUfq678
8IlKjPuIs8/jC03p+IOTs7OtBrAfZeVlLrQcld7cuwx2pppUhJGI3PO7/mKkasLsMkT0zQgb7HG5
X1vFLVc4SMh0V91Gl0oiMGLqamqwXQUfQnaPP7MglJAu+ateRwkbtkAetnyh8fn4/l89NC5jIQJr
akuX82BpDaciX6OXGv/VtYZKcnv3trVxk2+zS7xSBdJFizl4LggzUjdHGv48jljnZUwQDDXYH8Au
tIoa7V191qbNxTSd3zV44vl9dzanOXOiO23lY8qg82ZTjXeNQtCHJrcScEz7CdCn/QADCRxDbcXx
pRJLiOuYyiQv15wq0GNnwL2ihuVLI09T2P+UP/2PHKoHE0WAiyingdoy5ZkBfTrD/H6AXbh75QgC
eZ2EjubChnhKYRxTfg16sOhfK0PVhBsPwR6zjRhwX3VPJYxHn9rbgGYhWRGhxPBriyn33SWlJC2b
Jm6OW2lucUiO/ns/qc4flXOwDYD7f2qgxxErzWW9zOvkc07CTZQ45ODaeWj3uXExPZb5BSnQrQzQ
86KTu95vEO+6KZBFVaLSngypmZmpFwEoOeCTLbUNlVB8OtLed5C0+pnLbVDHS1aOzRKsf8V2o1pr
IbyhEOBrmfm57QZJjwFwemorEFHj1CvvB/zU7iQmuWq2Z5NPoZjvkR6xkD/lXHZePj4oEAcC1esr
O6eJRukiRL92JNwIoeX8pooQTSu9v4zu0y1h8Yvef7h/T3osSxqwr42zhf/J1rZ+tHG7xdCC0doH
e4ZsC88NAwIqybKccPS561qwYqH85HSNADwcC8T7bQK6/IUv5K/TU3Ih4PbkMFC4yUHzSsn3TthB
vC1jLdRlPf+1s1QPVXoWKIMiCXFvj/NcrJPtWg+dDoAK5ocWmWg7SB9PSpdnCOBCo0/5eW7J+muM
kBdRS11P+GsSghrNahbSVSq9NTuEJNoGzbH8H/OjIZc43jliUxAqGZfwtL2wUbtq3Dciz2+R92Gf
gx1jY/P2PuDy2oLsiBlHvPI3h3/9XStOsAMZ032efQYoJjfop3EXVq99m9CKChDQL3V0KieJWGf1
3I0RfdXWcsbcRAxNYedge30tZiHLWU5TKB/sc6gIqSBhdjRIkgHKI0EvYZCoFZwik873ETmz5s5F
mzXN6L0pwHvCLaUjztZ+BwKSDeENZAuUnLZbBOiMLSDvLhqqbTnDo0H7PKVfP1lfYgrTVwCbTkuo
6mqnLCzHp/nQfJ0E5Qk9CyDKwDnu9AS20oqiD4uYM+UjBvx9LRh6ZOzr8t0Z9si3lGIDCS1sNtpP
BO3Ewi9fOFryDNoo1a0IxZWo478tF4SBcKdwKxVND+/2CJq47se9WYqEkpY7EgtpQScOQAWKANgV
c7z+KyORrD3bFC+Qo2beJ3WFUZev3eHcSE2/PaACzdHv8gezH4DiXDEcvpmQ4v8eE3tTYx/i9PDz
SVrvTUkir0YU8xDBPAl8KZlHXvw/2weAYs9kprGJp8adT87p0+eievp21FCGjSBH8MfhR/LZyb9Y
sw83MZ12GIhbOCYEPPixds4o5v1bdhNhc0ehGevP/WOyvshnYFiB9Hgs/g9aecqE3ws62Jth8ecI
utikD6zE4XRzUxFOeR1Y5+d5qxxerw4x20jezpT/8BWrOW6aP6ujbP7VEVxLE35G96R4QkmvPU5E
Hu6tQHDsxRxZmIKrkkGUL7iemumfKguhuLcEBnnQWmGfBbeD55E3K3goxX0+aSMHP/3aYieIglkw
QFa6Eg8Yq56exWx4A3zktnSpt9yH0sYSXwk+MrLr1mdpDKEEGB1mzuZWs8J1+vkQXSsJm+sLDzdg
ATPz8954SGaO07fwDnyIeAuER/d/rOgNY1yitmWP/NOVtHL3epGsZ07Umh2APAfo49omUpaH3Ny2
Fvu7N+OzY8s7ury7FhuHDvGASGynJ+iGdXWaIx3h5jVpyYFYFYFQbcKH/o4DMb3biLzUsLiOKl86
Zfersp39UxE9I7luQLFIZwS0fzagCS5/n/F51GFe94ve9q4t+USKFBaoOByH9DclZSVBt43wHkJi
xIN7v75XvmmDYHT/cU4QfmKAMXB25XEIMlQO8mNqCk0bGdcfRhRySGjiC0yoNXk9Py6ZipaX8Dmy
O7cryAE4Amzmx1GCwl0Gkm/eN1+dP2M/Bkonh9LJiQYDHsNSa2Qy1OWZXOzduPOIvsgrvYdV7kfY
L4SlODxJDODctVD8yXqMsP8T/7m928UJ7fKQDSRjDQMxr3/NLDigbXoubyeLyujW20FBkOROlbu6
ugW3UR12B6S8Y52YPxD1r/bDSbYxz+96ysf2oEbdXJkP9CT1gOHbVwhXakwyfBMUhEk0ilh/WpUr
pmMtmWoDqSZ07M0dh3wwyhGAMiZ3v2m1LK7IyX/OWH/8PmFQJBcvPJuSpkxSGJfmtSdXJc2CCEnw
PVwC6gl2eIT/vZ0MI7hit3IpyV0K8/a0WzSeXo7a/+JfcJREDHuiNj2eHWjYGiDl6uu/PF6cE5xO
0u6K5yVr3TNIv0iGQGzX+KH+sAe3HiCkjFyhLlp3M0qqR3dTVHm44dnU0gvRH2V0m2AxAf7bzJDR
Zf3+39jWs7TuUz1y96CDxTHwL9JzCXJqWQrfH9KVTOxPjEgWjl2BHTeaas5YoINRP6GpP2NdDNYx
NsQ7GyK8BTrmRxi1KTsR/KhsEaoq6BA0WKt7Cf1kOAicAAEAQP/Y4Z/KhAGzh3ZbB7IPPTQi4b6t
6/IxZTQOIRWOy8qQ5koJIRdv2wTOS5wODLr/KI9SySyH3uuWCU0WKmjHJeEKVbjk8gPe6p1668Zk
ojuWI9JqJy9Vci7P+8hsi1D7jLjrPLQmx/L8x5hhatxeJ7BQqiO+IcCh9tsUpHTqRJqVb4DINMt1
eWNKqCE4VJbrcCcwy7iLRD/ZQPNMpZ7ny9OtXqsPeW8BWjFps+AyV5RsWBAXIRCgw36TwVV9IrtN
/NSzQYbbr+oHC1ih2pIF2sS2yWOGYQpmloeW65gCUAIpZZEMumryysW2xD+nmy4mGMhi8t63FACd
LIOha12KwDEznXss0+kaE2DEQVg3vQP5Sqvz/nXefIyqsNXEtNXqgc/Yizc0WebOHE9Vtt7vrfns
AqgmKCaoV7yq2zZTqomOBNEoV6YIvpQ8SLlzN3RKX6EOxqaXMdOQyQhFF+1zhn6nw6aL9w8phKWA
LnQbJgw4dc7f2FO44e8OMYxRGNWOp32HJKJ6jKO7gdf7DxNCMN1Riek25WSiV8gYNvAplgx7kzvp
BhplWkDMbRASFn23/XgfDV7sEtz3R9G0dhFQoM0V9PImoMtx2sk6Qh8z55457JYTvlixDFyDbGkx
jXRa+askDK9d6sNtWiAK/JGQ4hQuK8nJ4OQLhkTqVmuOPYeinJhKrHjx5C08p+Fm6YRL6amYsoOe
F9dlE6iUtowxPRD4XtOmJkz1kQ1p03UF9yL41/XnNdi+PSwZcCheYBIaY+YtjacLSk/lcRPhVabS
/UUTm6QHFBPTWprH0v18qlEb37wtnJGGMoypMJ3G5atJyAA2Z338u6I059bKPGN07ZLCl+3FM4mS
SyeMOLZZ3p8nNUjHpdp7cxAKy/49oqCFwRhuEYLGHYqV4KZbfQAYIlHCWQwiL9+5iVtHhSaHezS2
Ljx57W6YQEUWC+V6Kv8yapR6oyaZUZPcbi2GvHSMNNnzQO4pORBZHzo71nOV+b5vmmLOR0C3C5gH
0WzM0cxRu+Pp062qPidD+XLa8VTzt7lRfI1KI/hAmvoP7Dax7YruNPJPnrfbbppSTAaWmiYNhjur
dV6ukJT01X827Vr5xy+twefto9nRezIGQAgxbIJkAhQKhiAWGZcQDoukuLRdsdj3ozRTCYmtoILX
cKpKZnWuer7GID1/rrKUXapQF88pc06iTEarDrvTEwbI6VaeyqBlWZc0WmrjS9dsxitHFAMB5RE4
Z0SD1zbLKgR/9Jm3vEVXInLKYTG+1BBsV+HgsGMQ/SnbCIvkrA+TwiV/fi8iVj8Qdx3vt6b2C2rX
5KT1NzdnkL18zjHPOJ9Qpa1keMKYwAJMKKkCn6c4+BC20fBpOYeYNNTXJ8gsn4TFofjidiCLqtbb
MB8iLa+5zZZVszop0FuG0ZAT7k9IM7UAiu42u8Ojzf/3zFEE2XbhajN999Jht7FulbjnYRJOK6oI
OYamVCr9OGZYARgOlxQzqv+L25krDwJwz7MeekZ4XXceD0Aqa0sUkIv9Jvt32HVp6/nrSmD3DD30
LN7QJ3IAL82zxK0rXfiUSoFFslvVRBgXMRz7GK1GdFdM0gZQpOEpuQTwzXusxlGz/6rj4XPhkWxO
x92A+tHv+RWwM5OoTphEttM96cnhOSbJinxHoC9accGVr8l2nFttrq1H8vvWSODQuyRhx0nt6xts
tgrSxtFEVRJpMUFR5UuvQ1vTGjlE5Cix4Bv834W/HYho8VOg960dKx97C3ULDNf5G3mVpfZeZKUP
YJCskn8w8j+0I2/2QbdrOsjBAZCnqG0IWMByPDqP9G2G+a77aMjNAxMbReN+0NY9GQ3B9Y3GwVB2
4m7eVDUQ7BOLRNYBQfOgE9U5XQIV2VO/w33FLITzTAlTn77FyaTvLdJgayXagfazzcWL5UwExSZS
xeGbVd7AP1jKjrtaRqmnysQ5J/JZw/yPjlgG3XPg7ssmfpiR+jl1gIvZJw7dfkwLVJk1GSUMbuZ3
9TmoUdp/nAa+72ntZn/smJ7wYGvxvsN0c7kjNGuhsvwQlRTQM5yihG6eSOgZm3Hp9pLXSsV/qIVL
g82wMcpnvqLbjy8YGNVy0gWoq/bAq/xmtDIZ1wxdpbqYeEmm+O6eFdCi8yIotkdXXGecmINu5pC9
PUY/LgTwXps2sd4IuW/OaETbERTpp/Wh7HrXweauKEfifqC8onRVJGdQdGBEJg50KI6WHaslEDt6
1ig9szfc2WW+NnIL+mpEa0ryI104PNI+5kC8d6QBQhdPXDXJmgSJhIdJXg1AZ/19ScPI8f0Cc7Gv
QxLJLtOE2WSz3wPeMqU5yK9VGVSjQi2BQMYELTpH69nF0vb5ioK0R/WjqhNJ4jq8JTXt4Sz41mQ9
jHO6c8Cfmb3cSwi7SmXB/vX2lQ4krKLsG4QCzo0nXFFKxhNQwenDl3HxQJOQVp855lL2OJur1weB
oG1+7zE+nNOipQLwUdlnarJZ8xqN0odHIP70ciOPVuIxvR60OY5wuqr+sBXkdDYIfaCgtgm/wmKH
VwS7NXgPwjUpwTZ1iaFi9RWAwSzEanAgC93uDEnXvuyIkKgK6UgtwoLTorx37SvAD5oRFxVcifW8
qunLSXv/Z0wW3y7bREqb6+tiVFw+Vn7pIHTYVbLn0ZdGKnwDeo7o9kUSXPjRB9pn3AkOWbONTi/E
ZJwxWsLyQpmMbXmbXnNRICg9CqHwZ3Z8n5TFm94twuGKLEkvyPzqx0k+qeXh/Hbqsv87h4ep7q7Z
ut+gYyVfcXVtqZu0ZaxUSdqjiouNPv4ssbDVqt2ObvLkUkm+5f0EhTqzzlFwdoyEpzh5M8wmfGON
zlTOma4kBa49gQG+SmqG8GFwyTODpnjjJ/fsYruvQlePsZKGrjn/bXfnP/WGgU2VcXMuBXFvKol9
cev2gf7AGi4iYX+BtMZYsAaHrf4hw3A79EgGpMdzUSnDHhb5XGkKPZ1PhDbYLMH3YzeXPj0AvV+T
9e/LElYEyLfRKn1HIv5NFnzTFbli78BL57W3R51s3QoYARtLRhyeOLvYWSOhSgEMS+RJ5lyK9E2G
Osnlf/J9sTLBPy9n1XswqOckBtmFOH1KULIfw6DIYAdFtfYkfjLBVAkrEKAe1MOVI9IzYN6nT5lS
m+dEq9V5EBZ0dxSZ1pmVHTYwh0sWEVvu8F+VhPO8QfN570r/geMiF3ENPUAggn+M/4Q18n1J3LSu
+Oac/HsfNh/WAE7bJBVEyk3QNf0Yx7IYk7GOV9mo8MWii+hJf4DUawJufmhfzi+2kMcwTvjl3XLj
whcxUdrUHSxVag5VJp80dRm+igtuqdqV9HwPj/3B9XY3j8Rm092PJM4x6kKDJeHKrS0rKK4Rk2Qs
wnWj7NENXda3trLpNgfdTT0ILlawHwhp+c27h8viT4wuWsIR+fUWKRa5q5v+L9xMI8Kf/Lyqb/WN
g/vonTUa1Qvb2ZidiP+qjWwPL1NwR4Jpcfygvh0UN3b5p0/M/fQkbkAb0gbq/jeFWR9JpRbo753l
z9diFPoWofaKi0Q2HaG3BgHdUJPDQIM9sNPGWu1TQ87CKYqgGO3yPCOpsYEUcubU9QwPoqCnssQX
GQgzqKH2vf6jBCHWb5lHNbmPehtRqdNBMPgUmexdwum/OGjAH0saGzNJqGuketKqkRb6+hElLFgD
u7d/dFgpgxfbP/3sWKXPjGwOHUsE6m2VZpuDTnREgkJAabhaXkrChIN419fEfn/zt+F4rfQ88eje
3r4nSOIBQPMZKDW0r9nERInrk5gGpWRjacMHRgXAKftTaDfvKXhcEbTcT7hdJl87jO3qEAlfG/qi
oKfluUq/UHw3fpxE7OWJVnEsk1Oi6GXyvgfhsk3dIT8lNr35dvVcxY1SSwQZmnabJxuboAPCB5WA
6wupZpFw/yiPH7Tb8F4WbyKiDpc7D0Rq+xgtQsneGWI0n6LNPZqwrMbQoMVoAtZdC8Y6P6t2ZbaJ
1Ir+fzUToikHF8FbseNla99R9BQC8cl2KFUkOfvIxYK9CnEHsQ2NXnnu70Vj25W1urzXWM6vwVlK
dLURNqYs3SXV7Ri4SSPM68sqki6iOYoNUbTiujcQNEHOXHcWapRFZ7kamf1Yt2mjv9jPe3cgAqz+
cqGlsM4Z01GJjy825vmuybC8IJmt/kwJyjHE8cJcBdIejNkPxgzBPGnaXG4w7QXmeR/tI2c3ixCJ
pzutsNli949Hfce8tUITRan+1J9CzxLo7eyptpElukWJZ48f7LCwibahM8/+XruJiZAZ7ZW5U3nJ
B0eFi0u/Zc8zRkrue4tAMeDoPktyYvtWPdpShN9ZPKVqDflxbq3ykh49GMThdyv7rWtF66bgF91d
jKkJLskzLvuvS+jlnEzNUUOXasXrPvVRxjhOcjEDq6ErGdduIj7a3e0S+gypqZybe7lCjNIrSASO
ZIMIEKsP1rwZ5ByA1kZfYakmtzvSvTmpoT0ShQOG7MbtN3Eh/Ecc6ogqucnDNGN1BQ7MIFg4A540
siGc2W6fiBybbkytSmOsugQq4dCD1DwhMjRIK2u3Xj8KfAF1yBewUVtUGe6dkVifmC5UTauim8yj
v7Lok8v2+Am0p1Hr6qHNZuw/5Gr/JUUSgF/1ddODy3tDukSUZYCPTDUQZlktHXGDx++zw2/admI+
PNz8Nl8PgF5+by3tb5WDOmmbPYgmhRvPBITQW55w75tjE4fJN/IweejYlEi89QtA3Zh+OSvuDzj8
9gFraY9fH+8knP9HefGg0zzI8CL0vPPqvEKhvoVf6M5yHjBEww2rTsQaQUlmxsiYjrc/X921h4Fy
CL1SerFpQK0gP9U8kEX9cc+1ADaB6t4YbY/fdA/Q6lWF6mh/BrtWErLnp9dUvtdtcOocCaByTKXh
NvuFmr35cIfg5ACuDChn0WKo0Uk1EZ2TwjOy2grWxI5tfu9HnrjgRiJyG5c4KGdnK8UfuQadwoza
KO/lqFh5cEv/GiBpHSWBgzvUepbS9Db65oSgUSBDZzJ1YwS7mEXz+Grw3qut1CeQ0k3sSSe8jITE
+m1iJi8x+CnP4zTQQsbhx1NJnchxge3hUuaxUHoqQnD3ClRm90QSG8i3HNilih6tcr7TFsGtMBEQ
tOeYAgBfuoHXV0LcvPFzPPTAQiO8QtFCL0w4v12gE9/u6JSAwudBxJ572M9vUOOqJQwye1zUSbUq
2nJqWXPlASfiiazVpfYFDgNyOkL2I4ALhSanPlUeQghtULVvxWOzVs7/GNecKIFCo6EDn34UjWUh
3cJv2gwGKIAF0d0D9hCdayabjLllnQlLN0cHRHYLpFm+viBhHtgN46ECmQH8Nyk03XiCUljIV+nL
wgwAEWQm9f3rtXRpBh3QD1cYNbnf143Vffx+C05YDpeStNjyoEU/7AxajCLMLmqpJ6WqUb14Ql8a
qnsekTPTrdCKyxJQBGKIHrKiqy8ZiYP5+PwC56KcQySDcmvkO3iySjJUojghPJgmYiE56XKCZV6+
U3a3QGT4Kwo7vkO5pY5RjaeQHByRaSV9Jey2UkCqaHPSTMBtlO3aWzbDxYytl2DObhX4+hG7kijO
1T5r9ddA3Mi85xy2DyicAykiOFLx/RfXtQCvgfv/Yacs4LeB3T0bl7onMe8opGsRThdI/dhLu138
jwaYtLKctk/fCWH8vtn8Lm4Ac7FtUZrGw5mmEo9wIL4jlTGkgbXMNgYH057F0HuiviNCiVQn640y
iduBNYgdT9qNe20et5DjeFIHIRN7WdaNcelko6ZtDQJWjzjETJBOsZkjMZKtqCJyIhw4zbDvQR6B
g+VXKCznBeyZrAe65NPmtiq490c2AVpbuMitLnfazrjeaugV01sd9uRzrOoSqKURM+VUNU+nCVbV
TTYs+wVBzwrQntTkgR06ZsNPpaMHvc2kJZQ8dQjsEePNeuaPzGSf9PKd7WCImaDW1vk8I4MF/ANW
kE74lXf7ZjkdOuofHbk6i0bkHePCSRVcSzDJc3SGMs3KNwPyneH5mXkibaofqAyd2GdXVSfyarCe
FkqKfva9/IvyNd/0C8eWnMoRywUQ3QCUXQDyJzzplF2+VZtaQaNCjcoU3+xUjk/++f1CDzPNn8vm
9A3X6bkJEwlNo3dX4A5hmbrs6j4KTMBIzOaQKVDqH7YmvyZ4IeH36KUGg59P9LZmNiVU/BTXDIhf
qgk4B9Yla973nKKyQWcys+zLIG4Dbs0ofEggItttoWjE2u4k18Ttrsku9NlsEZFsMzg99JYcsySA
AkAKRwJIw/xAlp89dr6xKF0d+5505ATZzqDHJWNWjqBwjlOFO41bSSfCRif8srkqyl7Rsut6WuXd
7JtjIyiLjQxHmZKnsB3NdWBgbpl3TIIbdSquUtRCj9D1+JNWsemZHKf7hTIvBRwgUVNwjzf4Futq
ULk8bWUy55pIgMRmaibPDnvdvmQNuOwfWbOqOac6i61XmXF47RZTyBVB6K/oxDmOlnhCGOMDx8KZ
vOe3AZcsjHJNboIDRNXFf1SpmorGCUbdayMQ6oRJ9eHO9yf6kTJ4wuRtPGSb78T0YtAYEJMnSlxk
rTcSznC+wfbUqEB4VV7LXDLNmwhW4mp5+t4V8IliJM+7wO8hKU5l5WOnRdpo+VFbwdZetogKap+0
4jmIxwJLiURgkAQsmYT4fS4e4r+njZe4nH2REaaMEDOjrOli9PjmcxRa963uTX/+A/rrL0CLs3Iw
U1IqnUodgxwMgKqA5agDjg0FpHYGDhknH0kYUy+ze+aQpBhvu5EKKK/f4h0UC9bJTRZYis1+bHr2
+NKpzJfVEMw2u9l7etlwGXBbm00pmgU3FTchXismvNmw054W0Gf8qxbEk9/HlPYq+M7vN30CHeEF
qBN5VGTdWAO1pJgJcxl3bg7/dnTpAEUwq3yUHuP7UI0Mbb8Wcorgcr6H/JMovQfb9ilGD2DMEJIo
2+hOpaO9TyoQVnA77YeD6Uk62OqMKzjhkh8yYTTcjaIuaE2NxiSWFgvQPSMkN6TrSaNHqytTUPvM
8ZmgF18GW7YcgTKhKkA44B7Q1CKDheLmcwMND3R3VYxoChtquxT6oBEQvzNTJufv9SC9ejk3qGnU
UUxEtE6cQ/R68fsWcpIjnZkoFwmr8g2WYp8F90RV5nceBMv29hBI89VtE1wAUwFunR1aG5X5GAgk
jJREbNRKGLFI9NYyXJGwTkR696x4js/FQLOn3B7+3tDHjdo1XtpedKLpBhW8cSTkq+C6Z2jzfEpe
03K4dviYh0wRqU4qZaEQ/2kJAIAFJ99FpJMJn/wAq8ySwxhuBezmE8sjR7NixazBYfs5xV6AD8LL
DAaMhes8VfYN6eVaVYM94hMyR7fCXN+57EYVOg5FvLOvoN7e8dGLIopoBQQPwbj4n25hbhaboUmh
m/PYPhq2qbfYO8LmuK6Brfra8Zl3kEk50zWbLENT/e0GtXMWTiJwR2Httr28YPtSmpUDt28U7vOu
mvh2vHKf4+x4Oy1fGYgCTHBdQERgcaqO67x6gzPLL+8T+2LLPLf90e+2AazyoJpCaRCI7z6u1Y52
nloo2ENbbE7TRT+9v8IJ0PDLCi69my+aUOGxCMJM89luwsuFnjRSjKNik20Vl+ELisR7Yf/0ee/t
IL+gsgAslLX9DVZGhOwk2Uvsgsh6PqFtM9cHJypLXUZWTinBKLdHIsVlRQ7iNa3zPgriqaQMxRVf
DcSPgKmbnrYzTVneHl1KWjd4AG0F/MsMGc8+9B9SGQc1FZZOTtk5iqnWxHkmeb9PWx8Snlj4oQCe
1Xgbe4PXeIs/d8w3+2c+OnJz2VVsQ1DIOoFRUwMQgGQ96mp+7ueCjHFF+rbzbjrbyy5sHU24duru
CbwkjIgPPGy7Liv0kmfm/0u0wOHi1ELqyzD6lbxmAeGNcrd/p+JLMLUzOASqefaC0fPI9rxa/qBx
yVXjHLMB4TJdJKsAVGApfXE45yq1aVmK2FB8SefUg2lgHrm962HmJKm64ZusX7mVraegWIqvQ4xG
hfGML2O5E83IG110UvDSqZfQngQBoDiDXQF9+dFeriZw0DvXCsEAJdbkYuC/q+2/KVYCbfsjqHCC
GKirDHA2p3uKrMQus0zAMrqafnXNxwb6iYkysH9mucy8OtzGPAFGVNrCpds38b17j6TmC85imQAv
LR8rfvFrKcjlFuev4ETJeubTq57uvhKckDGxxye0ZXKE+P5xOVQmYpkxCmz5jSYXotNtdTLWThdn
vMqdu1Fo7ihWbGSteCMwYI57ZszgylDpglA/Gesebmyjf/GGSZ6pqeZETrg7qinFCK8ngvf2c2cc
Ls+WH4ztWwO+5xFkE6H9p5VaJUK1lwEANdkc6kmJvG8AhCSwMmQRzeP1qK+k0sa3gnFBkQ26yINj
FljUHvFGqIbiL/zxvAOrNgjfR1bgzsV0UyDVs4sQKdbbT+3Gn8FzD4Egk5eW72/qN8EhYeoVjcdW
QNSM7I7vyYBORba4jI4mdBi4qNlovOwkMq8jTILnGeEsprcWRX/S/a4LFxlVcoQss7Mfn7RZd1wz
jtIoUnN0+1VN0LFmvWxm66gLLFc17JxIB0mQiK2brfil+d19DqTLCZuntUSoULUj4my2oxVi0f6r
Owm61Q+g1vQU9RpQ0Zu+kZn+CdjZ/R59OOCSF4wv0XWD3Vnh3msVTd/s63PESC1bLLdlFLRPUavT
T4ZWMfNcrXYw4EOh6I6IXdcYAMjPZ280dWjs8OP7cTY8gs05YzHNS2ln1cMAmvRxWgCmzjAw/M2Z
7vS99UOU8Oji6wCUkHOBmsHdhBon+qlUMVHRagEHFRM0dRwj1xZDNHP/UNlxR4soY4mOnTmw/t/v
bjJrWf/xrW0aa/4OE3g+ncDGajiMCbPDei9jR6WQasd2mRbx3uGnvSUI2soJZIMkAMqREeOISMFw
6MXGA+0pNDsShMTGBdcl8bALhO5oUCY/CoLmOEO9FFO2U9hR9BLNh9NWLUAPbnOo5ztUq9XuREYE
FfbGiC3oMFrIyunL71019Eq3Qiu687Om5qAnJ84Gn64HS1w4a2+ZQB/8ZQAtPhjnFK0i3VGw/9nF
E1s+QOSxDYibYGDhgVQ9Jth1IkjWB7eabq6/3SHNvBZ1UOAm4kmxjvDSEGmyir/6mmHQZWe+K/Dz
JMhF/gj6LrChpvVDpnZQ3F7BwMuGcgwRi4Uawv2b3QKEAtEHzSHEYBj0KrF4gcL+pzgHK7/UrBXz
IRV8E3FCz67bhwscFLpTyJ06DbBcVBU2T9kr0VWr5PtdXEYErG6W+ptAYXRHGEnkMchtVhAA/e57
M1e27FmdyDamUzx1tBMuN2XY2BF2Ff4q2TNznx0YJ2sPRZvXLjIfQVJfhc7NAVHrZVdLvEa66xs2
qsbQSHWQp7BBuTpRbBrPFf4B4V0zr9bbBb9tYWMZKOU1iQFAZIHMzEHKZJzt2XN1jyl8S8m1Ul95
V55czEUvj9EZp6eR3JEjPkJmHlx5wyPmg2j/ocLSCaUy5iVBDfrZ/McrkmgYlr//NUDzagzzeIWg
9FG2Cy6YTBMD8VYqROyuXJhnKLLwRv93uUS2VIVnUC8gnE/kVFRMfK3un90Q+sLjBhiD+YQT4Zbq
Pq1HS/Ik3oWU9DABTe2zCTIdh9U5QyzsHE618z7dsxMXQg92oEBnp3OVJDfSHHGkPYcl0CNZqVLO
cwEmZSN5tKdUIpAO9layFCsjJ7kSa4ktAi101DYQ4DVwyVpgNrcBjMTEfQT5EgQ74UPYjkOW4+EE
SbsL74bcuD6RtfY1VGl+mGa01lKjmX6Cl7iyWUUt/vG6DvDmsBUCo6J2sJflPgAWfXhE0anxcAG+
yq0oDNZOQShidkGVi7QUtCP8NYyIs2vtPoXGcFu2a9rXpBktEPTIXrvEUeqlirwOJ9e+yRLjwXgj
PXkCj5nZOgjzx8yy4gRn0ULpO0Y6NFhmrs7ZRDgYnZrYFDFvR1nFOPcdseNSvnKR+qTATdg9hAnO
DSd1f34yXfYdgKM58oYKM9BEBQ6vHF91u8UblzPSROTZj5bk0TYk2q89TIEA81jCoOyjUWKF4ev6
KekVRgPTqeeu2fIfoqzAC47FmDilTmilFkrx4i8tw+RxdHPms3Eblt7FAbDBWrb3qivoD2Vcy6Fh
cBZGZSloP5dPDmL0SZzUdkmuTYE1NNiwyzG46pp/VJtIYfG2YxTr54djpK7BqYigy/NLXTzPKuHR
NBIMwt+Dxu71tglIlr9zVnQmrur4TJHwvOWA3WJybNWwYZtGpjuYRrS5bHieVP+xvVZeZrwtVxtC
iew2phH7ZUkANc1exBObqEWthbUA/TG3e+TD70g0M75ure0tmYQXyK84mSVpBhOyralzVVD6b9si
fxjpMtExHkYuM+CQ5lvaxCGa0T85cX2GC2mPwXtrnxtHlsGkEpWpB5tEFVsZCNHLSVU9kYOau5Wi
+fY2O2f6z7mltkYm3r7mNmX8q1f2KrYwtmr1PvNG4kLani8qhljAhVjNmBeIzJF+TWbD3DpQqKAL
pIEg3HNUvumxp7ya+voaA1c/F7WDEDJ76KtDkPlCrpy6hg78scyiLDp5zoHK9wiUKMdGfFOVRU3E
lM4p/jsFIwntj7CBv++cTCj3Yf2qerBz/f1CDfw3cXGvfPXZi+yOxShEUlnHy73Utj+w+WQTddQV
tT/WSpWIPRQQ1pyxq5vp0Ke0R7tTBcjnBM3/hN1gt+Mb6eARBjFf+YpgB6UAOze+lV7mXrRUkc73
l3iXdb9AknwWLqFBZILDo+e1+5+97PLGlIEyx6ejyK7om89G2PEfG3/M5N1O6q9gjuwXaspPeEVc
5ATXBiDWyTmtnD0aSALKt4pPrxcjV8iz78GGuaUVbyPp7XDT/NKztXO4vlG0Nb5bWYrYL+9iC8NB
Eb/sD2hQJAFdzlumIaON9NWXLtQlBh6qCLp+MoOPGKuBujeKYnNrcMih5WIjfDgoVgas04X2LgGG
1lsHI4knv5lPg5LWDkXY9Mxa748NV71DSwj5ba3JymtPGDiRk9Ozb3RFH2I/6Ap3XDjJHdQxUCEp
LuZuf1YidGF6mG7klNQZQ+55KJbeDaDbceKIetdhs0ZtWbSD15FBPJ/ZjDH/H74bg9jLo2sQVdII
qLeXoHHxVYdyUG/pNJgwZFZh2Rm7H2J65osTuJhTAc19UDOFnHto3S328pTcnYr1hPsgGBhfgtj4
t9SIcXd13tU6i1u3s3eQt6HApAzmd3xKFSeS56hG3hqUUHjNmF+SP1MprN7vwvRvD/aCUtn3r4O6
PHppBJURaZAvYSr9aVjy+JaK/8HJ1Mrv0Vka9/MFpy5kYaswssVlR5O0LwyzhNems+2u23B0+Epr
K3uzKbf0L9DdzTqNPGviJPHiJP+FX1sqBX6D/I7wqBziC+z9bJM4nWIkc95Uq0DptJNl/lPhrWWa
fstzNy85CG61JKd2reSM9m5XF1vqJ7Md5Id2ZEwIoto2SOPh2iIsFRrRbGVT26DftVWkJbmexFKV
qgfxXUJEyByUznYgGcz4oihCUBfN15A+dd0MBspwcFUNMs71BD1OPIcjkcw4LxhTOVLqjNzcYoeT
sw5j65Zs7wQThgyS9ekv9Lpud9AI84qyLi2oyp0A+g2JLepPExh8yX0M6RUWJxj6910KAYn1fowk
bdw8idShGXvjxDI7Ytf0I6k1ne2NkjOr355f0jKpjNsFB+vXf8q5W/xBcfBpnKpZQd3f2XtGTIa9
TyZOKRY2zlzM01Yi70PXPHL4jlDbIvbgb8AWj/jSXCxNtt3Oo5e11Zv3ATeNCjE8Gr17sWumJluV
kfmyYSt0ePP8QiJDRHo+hKa4jyRrLJGaM66aJOwNn3j/zg3w/GIBPnKbUrCCqFtbhla5XC3FzslJ
pP+9HqdGwkIv4tRsiXArciq7pBWWly9SR9sktNr8EI7teN4lpMMEtMGYGqrE1urYDEBv7jaWtbHO
MRBsTGtIi6nVspZfaWylCUi4KWhIlEblLj+gOt4RHB/mptVmuXwZ4c6kZMnv4RZIqu3TkoilZqTH
mUzCL9wR8LwWZ649G9K/qHADRHFM1wrhBzAoyUBnaIMGiuqPjV2qS6ez2mjeYRi/442j6UEbDZwE
t8PjnaSJmM9pjv+DvQ41ac8t1OdzwRmn4TMPj7uV46QnGXtFUr3MVrFmOqsuTp+VaDCEoBpmRxGl
ZuH/epoiLlEPT8UUjod1h9QezSUhZMELlW3Scl95SLusSSQ83v+wyaj1ItKXMB2jpZW43WBregzW
d4kDjg8KpUItN4EUWa7mcOhVj1oxFJ9GyfjtuViKarTgGkfDdPbhh076ucxevAFP3hRRpIGa9nDm
YuP3P4njwcw+SE2AP2n74Xn7gAopuLs+5PLHecicR07tqJakT2HuqTGS4h5wpzq5xHcfwwzDhaJH
gnPTes/g3xDykC70P8zn/zWj/0Onsvpc7kbeokx+O3qz+ZQBX75QLMPsgXZneyHHWa06qDeQnbXC
4ft6gOig7AzgRPOXW8bAJaKUXW5Xk2tTNqaVOpYPZGeBNQiaFYjSrgK5dLwcffajM6HDxASUqx1m
bnO1EOPX88KAl3HMe2odr46mhGJv7Iv8SczlNy3OJaxDCq5UG7QjpQb3AHmCoBa6Wbsr3xuWXqnC
3C3NNqC0Xd+UWPNsPTqK4gXlDiA7E+bBdDk1M3gnPvYOu4YJ3lLSTsQUAYg0u/Zo7o/XqkFh6LNg
4tlZ21zsaALJweAXIhnhwoloj8InlTRclZ7QUCieW/yNPlRoZh9C/b3pzM0xDzUUq7X+qz4n+cHJ
ezzSGzqyztGLZk5KyUYcVSVEQTKBd6Fa5X6Bbr/To2pfD6fx+F5YjCJakIaZpxmuSfssYA4GIQV2
tu5rbcKB95O5VlwK+STX3i+IGJsP3sAq3su/EDPB1EhsHelXlOxeVvtuzyi910ZA3sbZJyST6TXr
3j1a5OifNeiPnvX9kg4qccu8yUbBa/Cne+zlgJQrvyrIlm1USpYsZf0R+su80AuBcCDmuDJn1K15
aDjxUALWClHQ2wRy/pURznfEn+E+P5nzed2nKa9ucOF1ImLWkMeyIw4x22113Wa9gjX2ibjZ+9wZ
jNUzyiqCnCfXY5YKH6NHm0QPsRgFTvvRtojfRgosL+yTDAAivBD9XPwbmfhwV1PKZtLiSlZr8N1U
byoI7AwAfFrKHO2+DVZ10ZGnd6KcyQGjYltcfcsLcXTvvfRZ8CKdCSpO/ajzyPmF6viJtjlzHCP7
a3gTXogtFU4lf2g+i0TZFgw03r38ZVF+SwIcUZwOIAkc9p1/arYDBUVlskbHtycQ5StCHwmgkRMV
afSLKNofM87MN79700MRLrI8ifZYIUhF8b+yFmAJGoBYIJqbxTvR+2GnL0YmWlTdGTvTfdinOhDm
CaWJ/lYurjljOWT6vPUcG6DKjeC73N+lXtwHDm7HLFNGo2ox6OB9BQ4qTibp2LsXmk+mPOyIAEKP
YsIp4m+CbNkJ9tTwqsF1UHcEifezCueCxwyebqCsHpSXuN3qlkira3oWNeJONKTerUvQ15mG2+yt
sBulyXY/Qf0zXQhA5WUNgG0lcOIIx/oIsbE6W69xH4pzXESegahrMfbf9x4cguHw/IkddRSsCF4z
RfpyynZWxzgBVcdR50IG1wz+SH3+OSGUimWRuJTMocSd3jjg5NiI+P6ireIXWM8tLdLKBdhkYNEx
cfPwSnx6sCvB12DCr04dsn7G5djFMUPD0ZUrmAUQFBOZrfpDUA4bUzdGAibYLGT77x/3qAoCht6q
ZxcXhVEEsPgbkAxpzd37VppQyCPomv7Wa9Qf33jIgvBY0pGO7Eahm6OilJ7719etAuDSYhxiS8un
fTFDEXG7ion401Q8ccSjDA1ypsrg+J94LW74lH2u9rQTlsnm4qIsRmNw97pLUo+kQjfDdT4ovadj
+uSe01kDHl3RuVeNjfUrpqMdCl0CSvd316uPMsHdW6F6b5hkNzB6ytDv6x/wNtU+HfCaNLRWgZJz
/EaxVcv2C1Zwvf4x3hlsxe1exkmeql2NCvIpCMRgszoqTOoMBEHNAEorMjrIuUyQ8r1QSx8cl9fe
1T/w4tD7/eKTw1xo2+0Jioz8oKaVOnbsaRGZ7MW5DKfuM5RW7feQu7QolKDEvH0gE7RN4HNQKPjM
n8fShxsSHq2O3zGczb0Kh12t27ZuMAwYhuEWbHY7jwppiSnl3bUPsQzLvcFqmUG8LgIXirkk8HtM
zXneudQzicXfIqp59xaHWeXPLyMRA4yAzEfjL/astkj5IFPu4zQNnSZJLOy9OTBrXafLz2x9bgwp
2Pn9gt2+7IMy2x29WaUaQlkq0lrU7UeKY1DXtqMWsmmFebTrPxIOT05yBtNhCFo2UvWRrVBSeV8H
FxlzS8rTQesLJgdn/mc/SnckW/Y2i3/9qLVvSkdlvduHToHm+YFIg3vCs5V9gUzvUWgTOjdJMjxD
w4h9c6E50hivJrgRVmtD8VW2voIfgftOP3z9cUHjEyzYripY0TnoOlrVGA47dlLGtr2A2vqcuOKj
ClYZcZ7Mtdoh1t5NxqNQcB6+JpsZXcNlS/Zf6/lXpr6GtyBvcpRpBHSBPJjhPaDUtoukFKNWdFXz
BBivH97KlPZ9rQuPKaft/oEfvUZIEVnsTenhnLvGxhOk6hfTnfetXzqH3O0u5XQJH3y/DCz6bwSY
96belppEZCy0S88xZw65/32adLRiW9PV3yE7n9YRXoAZZ+yvDZdx3H85V/G5DsvjxMQ+URImQ4Dy
Im+kWP93Ve4Xm6vISEYuHN6YZBXxvc4SdAWonf8ehg4QFe6WROKjSmbCQOnhg4tsSvOJPNy3Zhl9
jkfV4RQKmP1jx7bhEg2HMmuQsEL/Vm2aEvyhMyOjeAOj/X07cZ7MPNGJqWsWc7nazg7FWvYThiHj
p/TQ9okPkrfsJfFCFRk0sm6xy/B30lBpvYogwdAHMz7dT27+VCHASNtGG1nxgWNoodm7DQASz3/p
m2GhGtMDMk0ugUeOWWTGhuGC9F2eWXZAKY0/imr4ilrji9M2WAx+yc/wj8amchVaRVVxCWz6LHnZ
E2dx8M8fQ2+7DhbGBpZSmV50mQjknbvB0+YErVU+J2UkPL/Qb6+eEVBMxeUM7jMS89AKx29A9jzr
GTGFsd2oNpykVQBvboyFjz9lw+3xZVb2G+7hTSn8U4n3UDxycXSw/hFhYjGJ1BQqeAPdt+gQKgjp
9lnKaH28k8OGAWLzY3t89dxJg9UqidOmGvAt05aSuEmqah1jTTl79aJiOmTGcfHbqK2m2e35dZZJ
6tkX3nkI/qDVVrRhuarqejVQccf6N2A0/m6JuRI9naeUrdP9ghNUa/TkxmAF2NsjrjqEeLbpLHgm
b2Mv4pVPVNEaDeM4yiw+TxUuWyoeU8WOqrRSo1pmF0cu106Lok3mgE/4PZUjIHeZquImOHrx5bHv
RR2FxbjsuKhjinf7A4ZD04rBncgG/sSQF99sOy/91DDuJB0g2pndF2PFrB2Z5+50/JQ3p7NHdWUG
Tx1AN4dZ4/7G91W8B08oS3LIuFB0/nsPysEd7eZg9riuST/oQTqjHSs1ztlLQcanWHTs1RD6BLW3
aecrRygixF6hJIkn8aGp4s3D3TLzoWIz9uhxPkWNRS3frvJmr4Fdsv+RUHNVFOLnKtcvy8vu0AFh
tsN1NkAO4Qe3eegHG3dpnCJrOBd82PmSSrE5nCvKUyFMdjCDi4iJr3zI4F46uj/zwLNhXarI0O4m
UHBEN04vdmHBRCJXYf6SOti6TgBxmgkmxcjUTi1raU7N/zM8rh239R5ZRDbcjJrZxZZ6yqh7fB+2
vdoEa0btuIqbZtJo6xZdBD5zgLvUWyNNmdkomizwNmsWTZ02VBwB6NyV8yjpAP8bSKrEN8rhSfIA
Biv6/Y43PKjHpKWoNwK5TuxPEmoYbKqzNE1hIsWm/ajLkDxdB9+q5STd9apv9qRV9Uw7T/HNUAL/
CSNkOXREuFod0qc0nPjiGTh77ToqiLO39U/yNqGRzBJrS50iM2o64crnRInbAw8x05ZRSMKTIbID
8ZlbPnYLp6K/5Q6WJxhgA+Jui/B4jtAiq7ANjvhZFwGj2VmQJHqfqbKQx8ywuBX0XmosP736D+3C
pw+JW8naxKbhiMYc1GNNCWBmj02KKfW8e/WcTeZpktMcMxMEw8YK/cg0nDrlgGTjJR4WzgMTGfa4
Il/NwQe/NCflcuYSfvAsS61cnUd1HPDCJUVB93ZT4Qmg6yDWPPDKvePwC3VkfpoXT8HRmvkO0PDF
tE++2d73zLVfMTbtjUcGQGDkCpijTVn9qgovUBZME0PgYzBT0TnEns4KJvEYkqlga+iI20V8vsw/
Bsa2zD+3ynaphv1MXwgiK0CzpsyorK9UEu+9RW5d/FAJGoZn68W4l/CCG9rgJGUlsfALK5G++oo2
Q68WJUbDTTC0bOd0uiWWlpkBKWYv46TvJS0Xe4pTrWpbK2KeqWAp8nL93lTjhLNUq7pzpDeQbkYR
GJtM3JCBhqwPlQmUo/066Y6lGoVTMfKZT0wJFSHjaWKp6PodK4BARVSBGyw9FjGgK1NS5v+hP1QI
H9VKR3Tm7t/fUTvvRvEyVoa0jzOc+MGGzKRRidX1HPwRE01PGcoGkrYbEDSlhK3MmLY1sNmeujdh
0x3aiqVj8oknmpqXhhKjzo7pVy27BhU3eoRJHuoMUlbDdJl52Ioryvi+2AThZL41DNWnme/lq9px
aKEwL7AHYhDq/xl613MLgFcKqzr3T4cndTWokEKMZnVJscgNzPy9ELUocA7FDfQObINot8BTI9vM
4Yju2nND6HSfCnVfEtmxRegv6k2M33U/nfMFB93EjRj6mv9dXQtfR2uwWrCUh9ZevJMgnufvLqn8
kQzYQchoQDNHKnWHjQ83fF52r9nxkrMnCFftB16sFQO1k8e9L7N1FDX7EXD4exj9IO71YGd/5lQi
Cq6lILXLa08+H0GukBbK8RCXeRkj41K8X86AbDLVLmWAPI8RsRGWg1EY4r5GqR6wmIm2Pwoj30S0
ibipCxwN+nKf+CEKUtZ28QQTZ3WqpUZ8HBwcZbaJ+k0sBaaf9Svo7jy8A6U4EaMCxki4NoTFJ+/9
kXlUhr524VaUimN1mEg+LaoIoA0ESUCYcoEeiSTXGq6c4fNkYrNkvWLAEQaVDeNXebFq/G2Sn2Zr
jesBBVEstT1yr3oIq/ZkTChRxh7OgkAbWv6YxdQ/H+ozrsrP+AcWKOSoIPG2bziSwziuLyweKZqW
nMtaXzEjHLVEyx/d3ETolTdHR392KbDlW1JLgdRS2NB7yqGVrkmM9oy+RX3gmIXq38JvBUInFfcN
qscc9F1Nq8Z7UaqgvbR79X0ZAko1n1hDpWOb88jPhMUAN0WnmgrHXEpMT0u2whVyo9TwgDxI8PNS
qiDGPiWmpW2AucEIFKS36J3g3NhlDvn9QrzR8EsUX2qZHf4Olo8ZSPiLj64KcuQPbnurfPeizFab
/DVDn028e/HKMB0TDc2ccC13FG4zzHAhg3lKna/GhEs6NtkWbqCSt2RF9ZvmlIOr9hNOXY90Mjrd
E0nDm+VthZt2M5wh7faDT9ZyE4yDxIScegTVLozgaHsM2GH9Gi5q2AFmx0w5xXEIHiFuF5B8Fkci
dfFO/q2l6Q73zNKqyBKIq6ckF6HodnM+Og9YX/VlJSMlaqKgVL609p2rprOwNEy0QwQd2WWh7DIS
NGLP3PywqUsEyvMbY4ZnaEKtMtx8tN73zwT8UsIUFVqYb62yB1pEHv+0AWlXqa0Y9cIijZB7DRQN
mjADYs7sAcG7rtbv9MAXVR7Oo4AeeKE4Sk2k+6UIRjls4sAKK5woU8yGNaWMltD3g6eX2uMUk14e
PsM99RsDYEyt/WcZATLqLJR7UBhxBrPpWPz46AqM96zy+i4E5wTJaJ/nE0VE4oKElL0XDOpX49U5
4cnVgiPwU0HHa1WnGHFCWivD14Nt+pWPJhdNa67q1+MO4hbfozIFiWzLsIUMr98e3CQsbZiAdXhy
3oCCEFIXMcECZh7la6SmZFh+WtvkMlAPa3kwH3GTx4OQtBKHGYoOOQ73MjYTlz/53GY5e6Q2KlDB
0TFLuf9BOBPJjkvFyQXpi+Ckm6QjgiZmRhhcnITkNJikOjnbSc5TEmNcqwGRZ7SKawVaz8rw2OIJ
LBwgNjJA+uBOt75DGLj9JPPrGLG+ogdNaR6HtZWjxrtBlxcAM6tJvEqJgL/CPKZ1MWP97TU8UFGR
XBjsNMcNI+iyKCSOQyRWLDQFPHA7s1rnBmhbUMAnBhZG6yRVHfx5sWCH/idCltQd/k14ZE/yofPP
BVCRcn/LPsuQHA63glXJeSg2hoEFKSNIC0D8wfFuWrj2en580Hgf/Jvm16Cx+n+7EiP8Hhz7XdRh
+JvbbqiwfJt9Gdt6WEwv/zN2G6CPPSYE124SlocvBdYW0egm/jaGrpKjmKPYogBrgJ95fMyQgbj5
d0RZQkze9rq/TfxWKI71I+jKM9G+DwNU0McLFOB5XZPjJ6bpW3qdSDAJfKtm1QTYhfg6rK9yf6Ie
aPDaqTera2WB06FGD8TL43IFByiGdk2JC8RBMuf6CtmFjYuAHAUhRgo6CAlpXzLMY5v11vGCZiZ9
HXwL0nixJ6je4HEKKbfxNZoP10WIqZ1eDhL/MzbQEwKGpVratdu/Xh1sgLWXoJMzfw8UTI2ysoRa
XvnbF14CNn6Sj/suff2g2ZLRM/YXjDTfZFwwkjaIY5DsIgPIK2WTNWmdaOm6s1mvKbrxs43J42/9
YwE1s3RIYtczT0+7FtHLbSejWA2rIlwQgx4qbpra2YC6D8/xeiuKmsOcBXBUovVvf5d/LCVLZz70
tsBSRBA2662ptOOnxP+2iQrHrarcT21yzOU5TkUF77Dnl9nb4bmZHQsa1eQhCRzZnWxZXm2ZRBXO
Ofm8NRFEzoRAN0qAClBPdGB3GkC46cV0Hg2UrRijoQMIhu2aOo/swse0oYyswFZT18tsMxB1oHdy
466a7a/m5YGuCLHqNCwsM/1EJHqlIw5oFIVD2yQkDXnxIdI6tgvmgtUmLqaomrM/6wMZPVfL3qQC
ZNe6PEfz5t3rH//9ncTqd1odv9J2cmqmH2nmkjEEAz89B7HWVks95e+JQlAxr/ZiH96+WOTrWzBx
03DdNPJZDiOhlMHKDdlUJcbSDhSwGK+FJuSwmrtu3xhb9unIMVSGpGbLRiGN/GjuuapU5mXcqIa5
/qlp6csoFRU7UU5fbuM1DtKxIPDVwj4NNvDO90uTYWUJcNVqGYVCFFDrYfkwsov6voPCRxPjirIR
qgQTuIuRqwbJLOZdPJylcucXbVujkV342D7KMbUOVJMYMcujV0hSahXkY1WZ3fQvG8IVA/P/7aBU
5o+F36sAc90SUjPZHQICXx5YI+HfbWYYtiUX6pbd5edJmkvMuykjJQqp8UumsKb6h430d2A9aY32
cAv7YYSArq96Lnr0IJlzD3X45jhF7ZUtJfc3H6QSi+9O4mGkoQtrwnmWC7HuBvD6b+XPIVOcw/53
zvEHaGod2QXCjFooUCXUSL+tZZiBg+na7ld6hZKf0eEaKGxIaeMU5A5wd/MZkYgr0w8a86kDcjwo
R8svRAussyJ/A2AdLyUAZyH5ZgQkYSb5T94XwWcP7qyN/sY2RmK3mYZLEkBO3VMakAy45wqA8W46
8OZO7ko8ICmxtTEMtSQaKrgHGwUPxf6ymVYhKWdPLut6NGefGBIQawhec3R1dOnenBnkurhPoWlk
+zryvUiU7sRgtcWB2Lx0PjdBAHUqOSTuYDPcwZXCFneV/hL+ryR4kK3Sezq5X7Zdk0Yfwd9KjxPv
/CxdwN+bbwL+ZYfU6bs2n80cR5G0rgMbTp+qs53nUl7Ga3o0F/7Wf+0gAv3KQfoETw6MPXmrEYHW
Z2/HCaA6BLmJaHbzCLGw9vGyd7fTWW32w8K0a7KuwsvbkzEKmG/r4BRP8pRwc1DIurxbPwL+56A/
3rvlcKJFRSB322cM6D7a4FJPGcYlvp3RTJMfCapTk5H2kHibamKJoBqOOAVfsc3U6BhjUObU30gk
3D3Hjn7Cwd6OYqsCgsUZpXrwa+EWfeOpZlxhYYAcq2vatBbM8wtH7Ji230+mZtTk429VAUl7yPND
aMFFZLt4YMdOKjibv2rI27d44UV8DemlD6zSxZ1pi1+aWuM2xaVYxLD5chB4+1wEbYlsfS8QznHV
nZZzFvvY4y2i2j6wp/YQzd03XtbgT3tMpt7+9QmlbrBsmz+v6hm+TvEg3ODMptSCwJX2tv998pKU
JgQqLjUEmrCkso1YMaIJLboqMsueI+AdUseLyWAaf87GbH1yDUNCt2XoMCkfIq8kKqvzbowhIw+U
FR4qvwR+6yEucB0zCYGqhSYFwQGdP4iYVp4yiyD55dPvAgABgDxXG+JsQG40GP2vkEjBPpM7FM9t
ymttR2vghwspjQvXikWr5RgkN8o+Tgcr8IxPXk9+x5rIZ7ezNKZS0mn4HsezPBbFpg+TxSOYKCKx
T1FtzI3yiAR/YTKCBsr+snCDX/hmo3t0GR33ZWX3EzOlIDsVfgmzi4pcJyV5WB8MqagoDum0HY1+
KZrS3S0RTVLHqsX/KFl8KMg8X0ThHKozlADox8XOm78aYMZ26F4hpCyEOXODdJ8gKTCgoEpF/weV
LEQ9EI+SPbUIeoh6jx2TiS3qKFhyrpryrPR5LgOFefPl9h6Vou/LCoRl+BTr1MwQDw9My07nPPWg
WKfWWuyHvdTFzmH5w5UI+b8IN0AUlYpqOMla/Eo4xRxbuVZeNnM6I1tTpasbVD/AsD17zOqtEii9
CTdHdOAJDlt+m/2GkS1QG5pr5QII8+mim0fAq6mWq+UT73eUTlFhlePWvw5yTH2FosnVcLvRsxGl
Ju4YpBIjQT9V610isGyfCTLjYIHCaK99DvTBTMs5j0k1psRiNmdqgVXtDPgdU1lCJTervpglgWi7
s18gehSjjV9LAXUASYyxhqLLdMZvPM0kUUpG6AE/l/MTWZ2oSKqZRMO6r3r55iZ9vVI7HkhDmB4Z
KgDhUqmHyIBVqezZiDemvn2oxKXuILZPNShZiCmxFBNjZhzlk6DiFcOEVj+QezB0OuvMpGw02US9
iXz0CWvFlTlQl9HWJSFnYchAU6kSXYsRyOSlWaEXKU9ogpOrReSy40hnu1c+n8VOUugQDP8PCIdu
2lMt3V2JRr6PUGmxHpqJICNeCRVMn7impqfrQu+ke/e24TGqxIeC2xLizMa4r0lci0Dyk6aKv+/4
fv+7be8hkcYAkuuYEDdG3SF9HcMlP3nPouScnHuyCQDT2aR+eMjZva4LpvulbwETnwx2pGdTeRFZ
7m3RXEcrciRrlHh2kTRBN5Z8txXW1iMNGR3K5Ivl29MCxCAmadFCuSYv0m9Ya1sZ2Bxpu0Ax7DtJ
3kILKKSIEHlNPyuIvJq8vylbCGKhzI24SUpUbv0slelUhnnF704rRMQDXG7zLyWdvMJle8ki4UTi
fnL2l7lCTro9NXDQ8V6wemIPOx5QJIr1fSZ3IiomZIr/DLWvx2Kq+6UR/41zRalbmfU2FHz5bRUL
/yqNdQzSL5cY+zQ01x6J6PHvqBDxu/3tlRm/6QvFFVFY1jw2Wcg+SAs//yYzuJDTAfOj7pttYIe6
EIKFSKH9gx7Uw9nPAzxot+AVOyqLiHM8Qlv0q+gJ4+WinY9mzwIwd7Mg17I1FZXulkJoooE+lnYC
I6FBt5XiiXWFX1XoNux24DWfJZEXZ7mcdgS3dDsbQKLjT/pIUellfhyMugWSSfGMFlJPOYaKWkzm
cRdMuNV2eWkJ5m26f0ZLCgWEJeghRotwfCD4UHfPPhBuwI3J0XdRdwAAMExmTqd0ahgX8piP8rDn
MRgX56D9D4fvUB+jCv1EeeFjgT+H7u1QvrIJ+PXabtTonHALSMHPnyuSyQPP4z9RJEP7dXJTMEtP
xaSmx1+YzkS9JopxGBaGYaI8la+m4vqCc2v1WTmw/xcpWhrFu9BbaUg4lGRO2MITTGuN/GzglwKN
RfzEUFvrd6P99kcduSOecTAfuBKs72hzpQ+A9e3ohXLfcJCfcZ2I+CvqAJ+Ce+SYMyr2995tMC2+
d1IBGY7nGG5B4jg3vSE6hZmzSn3B+HBli7dhNmiUjwqEMMpkfJvm7qUL0tTnzdbF1puyA+ejO8nI
86aAkYt6bFoNCFc4gzYe1DjjSQNxrd36d7TwUWSAVPu3+J5uPxw7NFITfvQZgFIlYpmp+v8OFxiN
y+o2zY8G6P9WncTTlFy14Bo0akCa4MLS0RK6yP+x1qjjvUnFZYaQ3rzJiSl8c82VsZq1sLwyUcS6
jY+l34X4O0Uhu6bZQtNFjU2C9hTiiGz30O+4tBynX9gHBjxfWKyPmNgop8mKuO6ASE5UznKgX92F
Jz15JNDHVqNyzXRF4wuHvS9ZrGaxiY9jSSKr/gSUoVPfXdhz6Ynu076rtXIjXUk8dT9hqPDLmvc4
GM7dZG5R1zUA4E751jobOOXsgBd0ijSjP0SJVIgCjns5Jn5Gs64+Ae7KqYxtfrylOQ9emOf6m4Ac
JUeoeclnOgcKHBl8HKrRlz/K95FVbmgrkYWAfLLNIwMWvbVnd2EKQjmHcchP8+2iZh7VtKwdgvSu
Ko28yy2ym+fyjBUBDvqJJHEidBRPxK+7euq2i3csMIqcFHjswKbVo1VFXceLiCb0lFbiyeLr1qfw
P4M2OY0HH3kEl2c9moQDYH6JB7F9QDCC/GU2eHrEGItAF/2BO0MbAfqiHC5omLx8w1wBEk4Ojl2X
R8iWeCxTwCX1wSBdBzJ1owO0KfAj4S5QVVOUaex3USzqJgL1k0K2cpS+cNREr5EBQ87eNL3f//qz
MytaFqwsCXbM2g8RLK5Fp+CH0tVOeDC2fruYKCtMP17CeBgYir4hEnwc1BbwRk5Ch2QDefnimLn1
0Hp6qhheHHxkSyX/fc+9k63l7jFsB51GTwqqJulhjwdv+E+S2dDXZp59Zgg/6pUu64p3XibBtlQz
6wvc6i/ZRu2u1Z2f0KKiH9VlwqQQdh3HMngnlytkDD+2pOA5T8J/BSa8Dva39DxS00SaIGQIsuV3
P5ejFsIiGzoLZM1tczHSJb2lsA1fTZcBi+VDLtmhcyP0Un0KcdWFR9FtoGMhBFsyFI+b0+IYcqzl
1iCT1c6H65BGYTY18uWYOlPI0hXzGadGBGNxZh1lh/jemHnflUJ/Tlzfa0qvGtFPh1pFdVWHlSwM
e8I66+8ITlEHYOcZNQoZWGWARqOfP/yje85p8xCMZSR9vDNSw052Hd6ENSKAj2X4fteehXl6L+Ol
gawMRh8uP/gKVWkCLnBavdkmqYm3NKOO2GHaPP0dZ9u9TTug9NfMInsAq3X6VZ3wyu3yfUvEjcu1
A5plWvywm4b9GESBbF5LbT02UySxl0KwkJk3UeLkFDdnrI9hDx02R/XKHHdG+2kSrlvik8wUfOfx
9cAo+TE0WvLcH9f/vZEcj6SZwNtqcc7gJa7dtjaiXmDa8WbMT3xXidIWepBY29ScofbhCu5h8IyS
cRksNRpUjSwEEHiDQidhFR9/TTl5glnJ2Ib1b8GRnlAXKe+t3Zzgm1nmhh02oUf7uWoZoBEczFKd
Aza4i49wPB7hEs8io3g15+PNt9dcbKsuV0eRZLP4nTQj2e6T/AXbSJlccXjxlKxG/NJxZMjxdILQ
zhhnVdfa62bk7+2pH1XW6/pTiayIi2rwDa0uF9Io3PFyNHCPvHGy/90sh+YZEL7AAKakuAytyza7
R9mqy5a+RsK4m14qvfygP1vBLy2jgYkKKLFB5666Zsxu80Wlz1sbQ0345ZL+TTrwmD3aaX++6m2f
Z0vNojbkeYQxAfeT988g84JsG/G08h8ZlmLOWKyhUS4fAZhHpBX89Ky6xXDm6qfmGVqzig3R3Vnk
z/++IKGrPfsku9deZqW0RNMCUT+/QoHoVGDauTIznrmw6NR2GDP5UBiZNuoX/CdD1LRIldIi8vPX
ca4eiTkkIjC1KB7Ju0vyqzkaKQQiv5+Mxr2JegVL3syAm3IIjjevtR0pmFXnRXfgT9ieHpgA47f0
ZSlkAxwg+h+AWYQ7E/bIzcVY1paXRn2W7wDnM8zFD/n/xq2szHYqbuSo6ETtRkrUFLHBkc4YXk3U
+B9TU+yIqNMe+xNsD5lMt9zbD8RcqfZz8I9iJZFtBLmlEHGkRFqnL40zevJeh961WHDCoPal4miG
7ZybQ7ke+txM70v8tUZTCicQaw2jTJ12JMomyxDtocpRL4gH/Bn1QEi1dakBAoLI2NIjK9vZCbB/
pARpP/Lkm3l6yEuNhuI2c9/2GJUO4/ZAiA8m8ihWUQWq7b/4fax+66Hs5Dkh1mNm9r1JTSHlVybG
tOTiSZTErCnXBZv/up+HAYnC7PWFTjssSh3CTGXGnpyxOlzMtzlTYQbZEha+30kfT1AgE9dNU86K
PB9+nPFtC+T8ie2fzKlYzx/jo33e8f5+FdxhgGQyHzJrIJQz5g0wcY0aerptaqlFZKVJb/T/6uQ7
nJUDIh5G2JQBDl3ZNj5J5lZ8MLvO4YoHl1TY36GGWSmP9J2l0RRgMtsXhdQzgwZ3ljUo1cl58XMy
bfSOJKDj5Toqk3pJ/vmQw/5c4w0g28s32VCr5piyvUq3yNpiiBe9huaZMVkywQXZtngT7/8ePo/p
xhaWvorzpdXOah+LS9iYmowqr554m7sqFNw78/Z16eeStOvc5Pchjk8tf1SWSRdtZlPaWvlOzOTR
zzV71rFNglNi9JX9vOCEyXWl1Gajd28ZEn4rKA1TTX46uZEAC/ieUoNLE7Ws7yLEP4i9BtAXt1KT
jvdk/j5567BZnjPkM4HM0gKeMbcUI3kuubvbRu4SeXWORwpyZ6jC2wozVtWnQCqjYxvD59ZE1OmJ
zAAWj/XoUAbR0I7gN0vr9rDWw68VsczsqOGG/6kK7zWO8McRkqBxkyhzUeX7UAaJ6a2n27r7seza
Qr5LajLy6cGA6zkEsVk6+UO/Skc76XDLGPVaseuZQWVCAyxs6ft8vAkbQQ1RL3UULyVK5Q65cFtC
RhVVeida6w7d0MxMswKNdYspLsfZji1QRGZH7xAZnaZb/NVtIG2j6Q4uehorz0UZ5/4cGwd7YvSf
+kPC+JCkER2+ZzR7f8MutasozoVnD0GlheB0Zy0MKweJ7lFwUXpzSf5XwAfYPWbtJr49IACrx0p6
j2fv+9kEbTueLU/V0JLfN5fx5zRFb9mnf+3oH9hKwRQ7jbhmHA7TLVWtjdDj0J/fmo+dxzvPrkVp
ekCczm7c0HGuawhhfLePdz9O1oS54smIVjJ4IYgVq3VJTnOV5py5BruNdoS2kxuV5v4VoR6yQviZ
lsN6TbKa9kb4vDLks7H79JrucUzT350rTJDputiFAEAxMPGF+DON+Rs04GCM0tw11ILqO9X+/qt2
mOd0ZL6NDCp3lLAz4ISC5Av9AzNuGWvIJ/bphHS70+ulwHHZGp3np5TBXKdJrbCljk+871MCB7RG
yc4LIFnPKfiGweIcp8Cx2+9CvBnkjoQ/IIN7nJmQYZzYF+kRnkp1WXgBPNF89FkEWvZxT+7a58PC
TVvMsJBUEUj57GdpNjXC4cBzURqKR0CTUwOQlLzlMXUtH+3JwQc3J3X33z2qCIa51UPdAdU5Fk09
3OqPIUXB0AQn2urGYK3RBunkF8yuzvzMkoiJ3/F3opi0SUXdMbZ+g7fl1StEPADffvLoreHSZbOr
XAnHL5DFhelysAX9iATJKYOk8IvXWNbvyhZ9eWUsrZXfRIdKF6Rd0TSGWXZEUSfArBMChbcpMnly
V6ZMMExj+pItizCZv6bsJQKXCH1Nb+gKwyfWLi9RM3MsWuOGZJsfM5TdIFU5va4OBasi537/064V
UjTP8cUZVnZsHGlqEMvrUl6PRFVog8nwhdxYDFvesWLATbh8Kci2wgc9fucNChnGtc9w4nIkY7Lk
lKNmTjl5bTJQgGRslJRPr18k4i7JEULUCN24px/DD+NxZ9/VQC+rUjqKhG2TVLGEdOrs2D9pQbVY
Gi0XkOg/A1uEy+Sm107vYA/htPEmQov87raVG/8F/3IZJvoQ2ITrAp9YW7Tx/drEXOlOx85yHIoh
o+d+0VnoyxOgsIsvRtASJnFtgd2/a0ZLA/FTF5SjVkM0mkh7eBQHvaT+Zgu92kHcMeoTN/wocVy0
k+gxExJVr9SfTz/uFm/cja16n4MstHw3RcElVDhDEErNtOYQkf8uol2j9fbYHGWjHd96Md5Hf4LQ
CBj1yYXczlmQEQmbJmlLI1GSxQd1WnxA3YNPkbnC9c2dvW2BfzA02Bzo9QN3S7x/rTdwg4VwDHbS
0GKCGI4fT7Nhe4gfRdTP6mJ1wLAE5MxAOJgRy7BAgZF/X4K+icA8KtlOGR6nJ2z6qK9lh4bubD05
gnEgQhY2CWzXN4DH+wKDW7twl8XsXszPx5tg+F4FkEP2fwWhxEb/34kQOC5sufloWSqun6Jh0/FY
P9w68WGFUMGj1Qg4scN63lDCHFNLtDmNCq1MDj4c8H5NWkzIBZyZbjUk2Sa1tVRPN4gQL7S2gifk
QWogco+IBydEraBj04JMlACt19cnZeR6qBKurRofJQGdGpGFjAYFQQQ+33KusOept/ZMUGdc4CH6
3Uq49EqN4cYc/gWt+ZvfsqvgiS9GmTpDsn24cX3dOrL1kOR4I/QdZgzY6spzJNZoSCR+0COI5By1
53CxINmxC3Gg8ubH6fBYzAVoGn+Akbp6FULuy/TYab+5y69L1wfh/GEAYbAS84TuA5lsWoglRsF+
OWAC8PjbdzzBk60G+fY9vqM+Etd46ErwsEEYHyi0g2PwNnrW4EpG2EiH058x2FI7ltt0ko4w1IpD
z5r8cMgQw2q8TaoCMwQyuajesX9AkRNMEjmi/a3euDRl7HPQ8vWbL/CdAgM8zx02VFP+mS78s0Hx
Q/mSR2amqNt6A2dOsNz/wFFCnoA3IONO0jzpnQd0lyqib0qiJ6fiNolju/u5dy3nbZaSnWOVyQj4
s8kqjx3ery2NWnt8A1jsoZgHEoJ5uYP5pS+Xmf5cvN9gZkv7BdcaV79aF+OxodXKCrP1uyewpHKq
9VhqjebVNJe6/Vvsu3VHpjyfXjpKZYdjd6c9YSO4xFPiia/bBHo/wJRDeznJXSq5WDabRKLjnYb4
8Ns1Q0iRBzMoZGLDeT1ZHGjmDVr8Aw7b17C3bc096s+CLcm6tdiUCIPLGjrI4wICbayjyD0UGRfi
yxBjqCTRzU+CSFCGptblhNn7KYc/JqEXxOvUH9Wc9vgmHjerRuGkYUKJvNDLOvtjM7c7ktxtRRJj
UFTKCUvZvFgBeqjCLy8abloOXUdZt9YQT/uLaPH9ToIH1/2ifvgx8xlsxom3lcAvHXR9AQsR1qmF
0ueHFKQIi8l9ls2wxkSnQqF66hSCdTXJUU0WwqkgXBaUKS1mng08ebwt+Y8xy76H3Sa0N8GwLypK
TLIorDCOSBg+YxLpo40IXseTIf/oP97tbFvik2bVsklOoM5YgSY7kfsPiKAs0gLMKODVeMjetVJ+
FfExxpbW9ZjALIwK7UKTv775VZBTHiW69uGoAs/sXmjLE8oXX4bsPB80CTJqioDDfRYlkPPDv262
3LqNI03azBshp8Z+9qPhY3qImAjxRzOUK+mhUwY6+7WGlQ/zFMQ9awQs2iKe8n4KVIpjlX6tHjpX
ZqWwzs+ObgUWDzeQVSaa9impEcxVahXI6ITnYkB3X0vLUdvMN165Jt9KAqj8kzo9lXVGzyM4sALX
ukpbZWdkeAzbgZ5kXT7YdiYeGQ2MAfHkn5NsxeVWPIZqUCZ8Oh/Fatu8AW0FwcGqCgn1ng3FjIZa
oZXXeDuiUfQ0Fdvj49ncR4BDMjwoop7Vs/yhhjFhWbDPVhpESOwbMCC4C4imLC4zkFDbnonJKJ7t
T9ZNI0PxlHFjFe6k2mnBG4x7Dvco9RUchqo33+Ck7XRot2fqCLsz6honUc15yx5KQeJ0rX9XoVxV
ICkWxiku5zwLBewxMHvQYNC+WobVd/61Y7uFIWQKkOi7lOPL+6AshAP6t2idHuFJLbh0X0aBGLy2
uDeUSby1exaMbl6BsPteJ9Xwx1MmwTl2nwPGjje4qtMnJJxIER2ejuExpeJAhHEsEaPFlLgSHB8p
nuKORXKEYuzP24pe81aw+zIlaZg+LnAAM2bCkrGSaCTuDEmzn5fQSjCydpRHBZXYBsoLYi30wrQJ
5Gad7G9b6ARiSlT2MkG1ynsenyxCHWqN1cuXiMvyyAjNJPqHb3IgxSIgrAP62YjiZNGaoKAXUqg2
paROfYIU2QHE7ie4eJ1fh4Id3hVIJAQMG9MGEiGQ7WS2ihFay8s/qk5afI3X4zLwN7GJEJivh8BC
xKRNkTgdnk2guSVcoKzpIec2cVzLndYWEBzbDerMkulfSOI4G22/pXsd/qFV0JRLzWDPWwgdkZwf
RtGfl3qkPM+aLvC7OJPH/8gvJ9K3F1JizAH5BU9etN4vTsIbnsJOG/Innw/19qzUwqk4kK+H+dz0
TPPeSZ9Fip/7eaWyfX2YWUXmwuqQfG0gdXyZQb+QqfmhMYp1m7D/ZutALwfhp773XQPDTxewcHFh
PFHlFGJcrgLeZC0RgmjUw1VVaHQ/mC8e4QQFw6/qiprXkX9OY2cGn7ztuoAIgOAaXuuYSKGWTZjZ
N2vexK6KE6PrjRustg079xGuUuIffV8xy7GxTXlPbc+bnw25NcY5SjxRuRDwAdUp97xPaZiFr1E6
CEKiaURdAPl6t+YArXnxqssbSdrByR9OVbz5jQ20r8rpKQ3089At+YKqE8QdSYexinggFSa1SMt7
UH5cuvgnerC1iL0VBROpF90YyP8dcKYL5GDNZ8Bd23NYIstHgz5kX94EaaZriK4OVAC4NrtS5aB6
44AoTSCmYqAxOAQ5HmARP6sU3HYuBmMS428ygiUf8zDluHOOPdXzQsliluxXYzkxoDw8NoLo3gAi
9VlTmB5qlbPiqwQsOZOFSG5aLmnjUX728ZSfhybud1JbZFSpAO3z3KZ7zEDlUA1HG7/SPHhFah2X
SzFnwEMun0NpRoM9dKtvcw/7Vdy/bGqOQbn+t2E7Mrs5ju8QaFcKCB0zCb2A1zaBHhcNA12BTQEQ
15ds1n8/7JzaixOV+y+xHp6aJt4NC6/vfEYwJgHZJeTCnc/AJbB+vUhWvMvgjvlJfcgYcojziMEG
P6hE5DWxKToNasoSFkqGzUXkbbZIYSHAgj51fo+XtJD2Ee7fjRouS7Ia9CzCjQvfwtN/mHH/fh62
TFGd84CzN+BdGXszMVQFC9s4x1UquhcZgFbXZTfvrwUG4vXdIDfT6WO0ZRGQmlgW60ZoJ9ZvoNGn
GzX8/e1wzW1vEIl4P8A/h28+2hWz1zeA9LeOBch+OlqxoVmOJGXqRlWFNBrUzjxbgmnWyLf3DMgM
FBFJ/S/fV1O253rAzaCzRFlNyFXQrnqvkH4V69HTBgtknvUFjChV6LaTTQ2O3UgZM060iATSTkqF
h1081hufjvoMZ76jLNf4VygVo4drncTDY3HR+hNrfNicZJgPHclNwsNu47k95RaP5WcegGHXz+MH
jIWC2+taLsdW4FfPR5O0XnIEG6RRZXlKVQkJz9TiwUeqbh3uruPBy/tu1nlKCnxj0OQ58E4/u8t6
WY4hBEGpSOVjV9WUg5R1pSJ1FKeq/3tOK/QlzYvLHkrfJJb/UBMVmXLTBNyyxO50rAK8NofqMGgS
H3JIxu2DxiOmkqp1bE5Ls7cQ+NfVojGTRCi7WWMrtXc9rwRnFE2RlnmJI2Dh8sT1tkxjy4HHMIuH
7x2H+f7uT+BVsiweiABBdMWLT1a8yQRWNkdICaKsi7C90vAS6vUqqp5dw3SbwsaHSbzqeGqNH8fY
CMJp40dFuqy61nXwPSub5zsZZgutPaGs04vMgXATPgRZR5n/7m4uhnNeHkksN1uFjYNkkyKWtCTs
DNc6otcP/JvrvPOvInOC/8TJ0RWPYKnlCZQ+l8rNYAfeoSJqnSOkILuVmzvSJIE9gNtssueqkj1C
stZEsbYCmF5lFAH4p0oB1oE6hZQLjQPVlow2xS2JAMJafqr8IW4Atm+PqEfG/KhKfFlbMYuakczz
fgDsf2gY1ItOxUnJgFzCeKjUF5nwLbjht1f4xjeKl9oFLYI2MR7T5aJJDw9asKbZVtoLqVj+KUYg
aqsGo96wotY6t88A9lZkruSVP/wmwivgVsS2FNCqMQ2P1D8yCcVYoumFlPzRksOwwuWBh9yxNza3
qP9+kT8/1fCFYoKhgXJToMOafIq2wUxnW5WwA9mSV0U0wFmvDAno7N0FDsQE/2GY1QFtnTphpsgH
sztOqneiEywqOlOtm1EONoggaLGfmedzULxXj9kxwsgk8A5ppBfkzcXNUKe3i1tYYKkKo+ZAaPjq
f86SNdLP62urVX9BYSbvIaK+GbhEzdb1Zgm9nRfeR9axBfOdLJLHU97GjPD3aojijKBUaI3ORBFt
2R8bnmJHma+iTH27F8JX0tzcJ6AtxIn/lWZhTMOPayP2uPgOkmjK3R4jd8w36bpFPB0c4/6uLISR
vrRh601KfSONeh8atGpsTxt49RRzTN0Bnw0bJ9ipKwfvX6oarDhUG318pfV7hKiSDQ4fSIFMTOIE
CMgVaqxn/0h031rEhNAYO0mUM4UVbs1YR9xIg73UuUAl3NAXw8ddJXBmOv77nhYJ99YcBeaeayRW
b0NjW8R+00lEUgk8yMZF6fv2wTKuLC0Z7UV0xlvxGejiVyJh6H/Ef7a/YLan68qWBWTVz1D9tsxW
if85yf4wI5Iuf2b6e6NmyZajxy3xEk6cns9DsSbVQ2bHNkwy5QDcFJM19z+2IYdpmpVhjij4gFyy
NWpG2tjMwhSp0tQYz5uTSMnEPeo1PaNkp5SG/KtVxMOu0TgzbM0S/t0qAt0pHVSeoNHBYpB2KlSy
nw8cZzS5HbpEITQQkX4UPFXRRr0igyh71SeNeJQfl3UeC7/jiZgMwCjm/90pjI5MF978mKDNraEW
KIKDjjaGCetv70g6FIubxB4BDEEBGsAATOU0nz2pwtp/JoySpaidDe/VREX4PstmLGze6tUf4jTa
yAdjib+zWPTuMeH2Q8pXji7uxuTkUueuRhUqAsz39Xi6j3ocwlm+y3Q+3VyFwKOp+utzJOS6lKUO
oYhwznzX4lyNTPWrL1T8iCxHBSEbbKDjGNF8UrBXyBa/hpCiyBswRUPN6Q4ObImP/B7JcKciJxMq
lNrom3bvkvpivWAckJ/2JjNENCKOlhNZROasHVg8zyP9x5pbsQ8iRD1ehPV5Ju+9b0ReK6YlRp3z
ECNld0Ngm0vukQBHsK9/HlDUYEwYMrRN+nXoAZO779jj1WekEnRKg6u4eWLVrBubbsu1Y6H61cGX
W2pgFoW/T0/949TNGY2iHjjOKBLP8WdrcOb8LQXyPTrHBxxHsUmE9YOei6AoyOBNNYGrBNjhfJ2S
Tt+F3Vyi3bRKdqymGVCF55KUFBZgZ1MO8kYIzBxfhaKTr9Twggk7ONsxWMKdlDVbnbOwhvP/C2J/
KXVDbmOQMgL6PQzRy7afRYuPaf4yRwDUP6xeBKCGO70aFndGYY2CgIcYP7s4tvnIBkEC1SGysR/x
h120HTUtZFwmVIdEHuinT5JBETsDYJhtDhVbghw5Ojr2224tqzDPtNCabU0JinzycOC+mM1sI1tt
xSbrz2zzaH+xWEkVBA/iF/qoFEEItHDpy2zlAznnhMBfWWxm3HiWzx6TrXrX1elJsqYb2s/i6Iov
CKXg/Yj2yKpK07utY/i6XHMuefNSEWDqriugwqQN+IuzaWGMQaCYYW3SLcgbadtF4nNZpBBilh5p
1lxQ5XogLGmUv+HzXPSulgwc5OLTKY3IN8SCrn14GAh+jUBDMyZ7u8O0JeDl8FAN7A+9lFkNl4FG
4eI6z4kClMUHmmt+D4DAhNW8bwqtgYZc8w9LgzCQq2TslxcK+FS77ZmoCujcJ88X8y7ijMzvE+C0
Dy/FAHiTFhbB2ppBcee3boqtCLKRYrt5y7dd+WDuVMjZ2ov33uTfNIMLnuRDn2j1LCffoQJK0rAj
0V/rZ1wF9a1bb0IVk3Eqa/0av/4ycxOzkRMdoYns8mRhJvHz2MWq2NwWuqf5h7Xg1jpzkcAsSQiT
7dfTfNww9kbQx/O700IRspcXV1EDAmzHGoaor0rdPUAzgM+eGJ4/EbaaHE27hfHqieY8UDUFoQyv
yVowMe07/fBvqYb/PVVsEOmO9jVtDbkVkYHj6IK6B3KjCyfsCFnwRh2MIVvy5gE6BBNqmhekE9hR
bqnrCIqcCFjJDrJ9Pr9uhFWJARyw3LdIWtWXJc2KGmcd83je67pv4w8ooAfFIx+BgJ32dr1LFICN
kSotNNhKmdlIY/tG0fVdSoswjjM6qy7QHntZqTkHAtNQJ3Sgibtsfm2oy+yevDNnVypKfYO27lwt
Vk3ZhOzKw8a2uDF1SdLeuyMseWE0QMgwFbYNWAUP3Are7dz0RYff1NHvxyepvlWSVF12SmZbyS7U
wMELhm7enJHZUqsGyJ4t0N4kBRWdYcJKLE72vcULCFJ/Ha1hGi2szF4sDkzJ1y8OWm2VfnMVq7J+
AgsNF86Ev1vtC5It81tqRfBVhTv+5w5h7J1I7hlhj9PBefQdsrzzqqtm/SlRpNmIn+/w6F/vW9O1
Pi2G9FcEPRwZfyLH0o9hAqDMYN3zVuHcwjpYB620Fjo7Yz051IoeKvozgGcCp7dVYM+HpsAv/r54
qK1TLr1MyfVqAgqyl0usLtOvGBD36nG1X0jzpHndwfyh6pVoAhiyOycxXI04LpTOKd+N43vqOHUR
ejFEyL0FbThLaNN4EM2wr/DX6U7DhZnzx4Rsf8FxIwbHvFl19woDLLgA7zqDCXnCiU27yBsGjKK2
arKUtI32Zp1e2Gawn6GKZL1CYgODCnf7u/Yita/IFoZwmEtzyi4GRZRvWa1Y+rdDpPkLCeEVuFn3
1BZhF4Q32Y1zSd2oDr+uHx+Y2KaZxp2dW8WWP2elzn7RNPn9yrcguM6Ft2sYIEELSwj5jeWiwxjV
jZMJ2f9oRSDVy2n/bEOmfD5fnUVw0gjPRXPaA/ZSHWrUw3X+DdUCoB2ntQmBbWmpotzzl7J3JLwg
sR6SZzc/Sk8iiGSrhKDkPynuRD68gtRqyjocg8/MsqIJ98RmxpnIit5fewfHfwgA+XQFLMQXY2RO
SlNt9PSPjWUcCAcaoJk8+gWRBNEdAgsKHsjHoTEizUkOIeUh4wzuyi/lvVQJp0TyhCPxTGT/c6gn
uI4BOudJtI+iJeVKSYhwHvuHyEsJG86Vq8sp4EkQ4ILKiAOO3D4/OoL0WQaA0uagqpWLC7gITbpp
B634PlPaJ+Hw4H/56pdCe6Y2D5/iztOYzBbSRwMO+8aHkmZ6Pz/5dnpL3FzedDogrl+C1iNf5qxq
gMgfRyRKTctdNf6GiXYf5Ffj+8hkiv3bje+oN2yYYvvCPJlevf9mi1XPClaQwen9ihyOBU5lU6yp
PDCIDGRanGe8F0u6vPiQRHvWg4P5o2nbi81P1AYevOpgwoMwyEepC/4WwjWQjPvkgk/Kj6Ztfhsw
ie6nzBGEMEOqRzdrvDfiy6tykUdzGD4hzbcLDAP0aEqiFPQ5teG9HPy5ck/efHyqdVzyb4zdtDsy
SmZf8k0kQAxbxzVHESyE3rzabbx+q4HsNpElkKYIYCEgwbo9pfr/T8FAy/WzpQY0BdR97ggS7RXq
xYGdF0VH7XASj2iH+GUopWo8MHTo/Q61gEmPkbqYyVHA0/oD5Dj91OZZY+SGK4wyG8qa5ALAyo4/
8vQXpP69CHxw8He5GKd2/V6AjHzIQ8dVbbByI3RH455paHNYzyti0yLgztG+N+ei12i5HVFp4WqC
N9WyGpCWYq85Q52rHg1L+gRWf8sbxCcit3eaoyqCpMq2RtUypTmBjMwKRRdxKx6Ynsfkum1+NI1I
UHoZwDuzYRJOQ8NAAw821i5h8HjU94YIYeT1F/VrmJI5zgKJ2bpHZSf27kEXi5u8tBhFIDLX/HXB
VY1/z+b0DXeOUB5kDby6gvJVZL3VBEND19BaaepbqC4ew2nG/BOFHkA6XE8wdvSD5d43aAtH1Fk2
DiCkyYxw+TVb/GttiDzGii1jsXCVAunCi5xZzdXFkgdsxdjM9tNONyy1fqLVsOZ9HLSML37KkVju
/PmgjSKvH/C/IAB8pz2LGNM/Rvs1iXXEQTST10N6ybvd9CXcxiu6Sz6lusaBMv6rZWzEH7BHcb2M
GLVVyiPv5OcUZj9kofBU15lcezmpUyWhmcE7DOd9jZwunJ+ini0mLVoz6Zc3CMuXWTWfGLJcM1jb
131xJNKlcoob6QzsZqf2AFNE/4LtCHdDmHYNFReusbb9+L8/XMqVQa0qKQaxiO6K6hF1e8/RuP1z
n1To1tceQPxpXRGHUi6P7bz665fHXf/nunTVbCEvTaTE54z13EPE7a1VIK8ETBLU5yWbumS3CDi8
vzPFixjfm71nicK7wxSxJAOhdEOnh+v2XD+3J8YhSnxxdoNwGxCV+8TA/xrBarSlgztZsXBNzUxj
6p2EbQkhC/akLHw6n6HsSFgQtCwz39iraWuTmrL9pjBQdqb9VAnd/nw/uwtpli1IGQXF71Q5cLi9
aollHq47f650zG8Qezq4Bw+DCFKBwWu/WROxHoy0IuoZAeWxRlI9LCthETK4nkKtlrXcLbHkOvQk
+m2yPpMKSWPbQyAN/TnxVAOeETbhOrkcMVfl5AoHXsebkrHK8xXAe5TL90pTra98jmAd8flbU6hH
k9g6bGZtLF/ahQWYA9zsgpBtV06vZN1tmZ77R3cQiG6oc1OzmzrgZKc2Es4bRsNiPfKljSfrFBmw
Q0W59a2xYZjvVKGdaJY6VjEufiSTclMjuUjc43I4qHCMW7GIfjJ3zEXAIzjN7mWW4GhkKGByoqfq
v7son165pk5drvwztXjoNpyYqECnUvoLaR7co7cwUwu0e89dkGU/eP2kIU9WR4FLxTS0tGyMv52d
sY8M/uFLw6p+PC8Rag8nJeRIGxxNJUKqY4wx80bJWR6AMKez6KVVLtPNWWY82gJw5j3+Vn6vACVt
H8Sw4DWjmnCsWxa/gwOy5k48qnNeWh6D01mcfCu4N3ZpWuaO2Yr1/pe1TGA1gjy+X80si/+JaDBl
AsJKNCVP74kR8b573eIehtoFgQIVEMACFUyLStU20xbyqaQVzIyC0ByeIYIIeoq+xIyUp6SxBF3/
hmNnbR5Q2AHqW1/Rn75Bj+4dQiDXActYAlBQcrWGPYTQaNmT2EnbRD60DXuD+NQ76NVa1Zh6S1gK
2624cVJRVHU/NWbXe9EmlD4Qq9gGgb9u1AA+XeQcfr49NhNyuaDwc7TUMRDXP9F9IFNcs2lGGCAq
cNJjM6OkZFlV2ipdRyjToPCF2GHfLGXEdTGkmYS/K0wgWKLwJv85BgYJoDioM3qI9gLl5HFSEjoE
4nAhYLC7NMqXnxRIGHZLWby6v/z+yAN5wFCdn0nKL6xdy05ygghaQVI2NWRBxHn3szLV//0mFTRD
p6oOw11wLpwZKZ3LutIskPj6HjcO8PZTaUkzci7qXaOm0arkMzKgxZNwVnrRlwJ0cgxBmE/4ddV9
b72MRTb3z0Nil5wZuS57qqJF1gF0QMjNY2P8flZeiA74GiUcbbVQDNjqkfFO+Auvr2FLdrlpjlv5
W1jaUhpobE91NqaXhduug315dAZGUxQrlMgQ3o91hDxes5W8tDvH4sB0UnQg+m8ZcnEhAZ7qOAJu
lnZAORTxNavCIAhBWCD5hCoiGAylJm2yxwE2u9L0guCOv0wRQ8hMZu/8igJqb4Ma6tmplrNYQW5r
wHSX6azNmkXNqQhIhVbUV3Bz7cMwlxnstdQXXEhrgHptO9joVxhrnZHB5U+UPOv1GrBcOkQ1BxF1
1n0FlhakKN+Rf25fj7nS1cPWEtdp9hbR69rO7+/JIK8V+Do/KCgjyAPswFpxYTnd8BOMVuGmlQqp
ohMHhSksjVDHX7fCa0iWcQacQ+q2EE9Xg0QF4nTJdwNgzR5wAcZ5hoLxcqxNxuV5RUrkGed5NZ5q
SA8nSi+skZPgoVC3tBRWJAilNQUxYebwpxjqmOJHl6zc3P4jZygjTwTvL/A9CQ4P+wbi6umyVKL6
vG4qmPfQ/aEU1+wBCCfJhHEJR+lexTSSADxJppSZfu0uDWhdkwq/bYN5a79Rl7WZFoU/DvDFeeVB
jclEuuOYPrQx83AlbBBakvoO+gEnrCW9C6F72NFujcXHM97cp0iwUCSS+shBIeNBaZwrpm4xH7wl
dy9XyE2cvz58q3HikwlN8/T4A84JSk4Twu3qs4qCLt/VmndGKCsryASIzSgZ2cMMBGhrWtHANMPI
k3P+8ckvCfWcvmWUzG4vGnIzVD/jaG5AbDLWkmUpDx1gtm1++LBKa+qOd94OboYFvsYcScTKFzAI
zLGuxTasYS2LNdUI0cvdxVhSvgvQaZIJdH9fWMBWNtY8++1/XVfgEZrEbtho8VB6azz7YuPp9MK2
48e2FIFqXeHBJ1TxmVD3KpYb2Dr5SIFBgoB22qCYf7a9a4/MLDIJbzHf7u4rtABSWQLA1hAYynO1
n3jZsb8656t7TB8WzJdeOLjfz9L/ys8rTVo2KSCqzXq1XzNwBhaSEOZ2Vc1rTXUEAjNXpDqsqWvn
eRL2fcb5RvY4BuPB/fXYNf26gfXC7UQWQyzaQG7GC6w93wsVliz9l7bzyi+wuhfak9IyhtnIR12t
bMkXdQ7fvPDxXFmZKAyDK4w+g6G7y3E8Y52VkC6kQz4NxsPfTXx1Kq7jyy9bD4vgTmk4+AEWvMvz
LeEd9hLPJEBOc/9uO8Ms3PQBHCfjLdWeNKk2VX7ezpU8WbZqjujg3BPWE6XU2MVUlKtgBe1Glrsc
cTH5YzhmEImC/h0xxl7SkigssUDTgzi02+TSJHs/A09PcFXkvLGZC8qHt5rz7tsNaUcolj4OXvHd
ZUuEiAP9tFpgwVvzwFNGf826SPFGYYc8PHeEAWhdqPaBu6KStL1K00hKp0eHVZbIy/G4TC2VPNxI
Ro9tjzMwFZPss2LihfGmAe0wQBbBfydFprrD5sId5JgTbvo21dDkbYproYMlo3g1WJ6QJSrFftv7
mg/fa1l0R5xyRBkOAf5gb5w21jQJAobQfw06C2GVY69kdH+zdfoYBIJgd59DTw304XRpaOO/VWyo
lMSfK/s63pwSg6WIcPlKwuW58QeINXZBRh9ZouG1lW2oDlFebz1DrL+iqb3KjOLsIiB3fN8urd8F
8CIP1Xb4WJQiutk4nDve0pAG1aZ9w7+tnYWBiEe78WE15C3BoV012RYS2v/raX+0LI8pSrb9qTaj
znuPUiowBO/ACY8kEuNgJ6YsYcOWg0AUT0OotCG8mLgG+WjfIh8VStK7+U1CuHLnZJWS4qke60KW
eYCo7Fw1Hh1QSjeNam+/P0a9FMPggrBjGtx3yEwoEioygiZrVR4ny2YQZXjx/iKbbwJf57TQOqFk
yEgWzYpcdz8mcMb8ODzBmpMFoyDJLsFcZZ33xU6X4AmEG2bNNp4Y67Ez1+t1rSVeAbf1nj2wIL36
rVH2J3MxWeSaCGIK8Qn9fN5pFTtTV0b8Dj79TUsDDGgomGkO07itOJc+Fjj5KOz3Oz/YFBlU/ual
Se0/vvJVZkOscJDIgxDZv6CNaGe5JhY2417Gla4dkxrtc2CX7RgUxXvP998FOqKZdsTwWYV94IHY
neiHAu8Voctpj9G626ydLyNdG4DEYgdYrLxzQJqtm4VOdkMGsByfGqz8iXyVWzX4giK7sghGv1l6
wUJVPwAiwcE8oLjJLO62dboI1pNgs8+p31RJ++4brcQH7NgZjSsktjyYp93T6H8TBNZSFGRZGGKT
7Z5Aig+vHGxjeUYyS6oOSbyfeKA6nVgksOgmtItyzf9vovMh41kecWDKpd0woIAu6G+tiWwjNUtk
BfjNlV47M+9hrHbUpXW34GIagYF0mgfWDKHshyU2oC4opN7PLtToH2fQaFokOL0b8QVgk+q9LYlH
N7/ETqgsonfhfK5F86+wl2nvC6rZ/zQeqdplxCTRfxc33bYKevbUK68Wrud8Uh+YL0fsd7cdpyWt
HZPCgyLeY7RMo0oJ3UhYssl6eh3IaAaTUy5Dy12fbiULcF7OqSkXcRvgvfe9sFCrEOslvEFmJy3s
RW2wNVHxZ3owhhBQ/Q2bUSuPNtg3Ptr8UEXzWe/P1ycM6HnVL3RwuU4//LzOLAMV8XTWoA2bteXi
+SZ2uu/jaihChdFArKrFDuyP0rP7rmlWwhZv+9LtL3fQqepLH18I4i5CVLw3Q4ux6vnTJKq0NALW
map4034wmUQx5Y+pU5oFEEKGpU0w1vb4RXWkuYjOQalwXqyLQlqaBDD9wipZEVHjtCtqjdFEjE+1
1uZZxSv6aGdO2QKVvNwlBgsZkk11TzPwEa9yaqkwLNOEB1uMsPFZaCx2d2T1ON2bkPux3ldsnO4H
hNmI5eZes76++wdAaxQU+EC4wUzO4OAqztPgFO+YVxn9umwj0gSDQFw1sb9tI7R/NcWwNUrTsP0n
aMqkeQ+6R7sGuoRu3p/NJrsxUJgbLljIODxRnWzliky01S6LKAfQ5GPSjbmGY9h1Yy6pIkGghhYV
Clnt56FgYAX3S8pK1YOwxw7YLhbIEM6B20yQMVKLH0rJf7CGJPbgnjfovPLkfh/5JvSLtNfw8Q0E
1oX7Rp/mNxHO8wxCOr/7YVIsTePXM1paRChVx0gjdYhax+C4KO8VpmxsAn3gmDDRkhOMpbHui/Eh
2yS5wGVOBkRMfHzB9rnsRZCNH7S8cBvudSAPNlxJBa1qoCCxVjK3mDQZH0FmEXOAlZ2+SeheqBqU
UCiXBYKfUU4tAyzxoB5BHUAtW7C/d0IW9bnXWDgtEiEhYweHrdalmVDqNRggpoiVMCqmIr8gKPlG
pWIpay0SESjiNs1wrIr49BD4msVCcSyz54MLEIWOuzeG0AWeud8a2ZXI2l0/q+bRD88Y/O6TUia6
AfzELMfMRvLtRBAHxk2DETtrxCSQlwXGchE25zzsHXlW79OVCkh7h9bC7DhhLf+iEU02DyWgMxDN
bLOl5+Bh/fzOWFMmb9avpCaW79o755iA80y0jSkytIiNVXmKhMdw8evz7dytn0vMxtfVRQMFyU0D
P7pYVpsePFhD2xFPA7nNKqIBjaVIA7XjJwV0jN7m8V7evkka05EKVb6vzufX+/sgC6xvrFhc+ZEf
g9yV0EMGPhhtzomN1HPGPim2b/adbWm3Leizk6wwve0o7vWXQhr7UNR+4vRcdfj1+I5AgAvrgp89
4iQsrObX4NoqOOIuGgZmwRzKhcCzUSowentlqAuG/DGbfNtY3QFmJEG++k+Ay6hMtHxrW+RKZ0HK
wK3c4qGAsWsI4irePnvlWWVbBz0XIf6GkZ2Te2OtYyreQA7wlVRvepwCGZYhw4fmNVraKOK4fK88
hs6k7Df2O2aNbjo+DSfunBA5Y7WUqg2kMSU/vGH3E/RAIFBVyzpPspECqdZ3Z//VM9GO8Nspie1+
Hldxnab/sdL16TbtYYXVbIUzh2T8hLdwxz3WUKFB4skmbvupRFuuVTCtCNoABs2oK2znb/AubGgH
Frw1GiOYzs6E6doBrE6HQvicZ9pC3w2Nn5vLzGL3BnFL8xhcfuGsqNimWTCAEUWbwot4BdjNrKTE
REGjwLzgD0Rutq4THo9VfOM5s3uoiiMpoQmsENHbohlmjhTVQnhvKeAcnqpR3zuaOQRnz5YPkCjZ
Qx79l7hQv7ydwUMGBzmB7vIVGxpMuiR/2ME/9gDA8rbvxfG00ILpfzmVaxbTDfaSiQw7pJeAyk9u
0Kd41C6ucggDK/gbO4OBsv2+JWMl9g3MEpfYyvUxQkz/dAXsujZ2SagM15BwXcnzJnqxCNQlGe0F
kSXeNz5pHmwUh7lX7cLfyuyLXm2sI+7+P/T/IWCcqiqj0y1IfnrtS2GbG6MqVXCZc3vW3ZxL1fDJ
Q8wMyDc4UyK/+hscR/RYBhMZKmoXN4MwI0+d50eRcvtd7dTkGvDTN+dDCpcarNVfweyOOwku0EvP
BamDcBGr7fnIyklXBjqOMoqvjSvJyvraavQHGm7HTeTLUjq7S1kfrDTePoGKMszcl4fKJ2AzJWAs
AZQblr3f/qUaSkR4pYQl/zZCGnySFD9j3qx0XKUhHLImCPvh4YrEj0liOdlq91SHPWgu3qG1IiIE
OeD1qjjTmkkasqhi4KL16rjaJznrwjh4uV6L46LBkn+tdoDxKfjn37rrxzdtDW2YUcYptVcXQ5U5
aIkWgQnhlOLRLVv5PcLlQdSWlOmI/HFXENMrPy/lJYL62PWeFtT08U6U3wOhndOeVlXC3nGG5VlB
5Wqc5kKTOSDyAgDpoRmbbE3KXO6I+MGtCMCitwLMqePZJMSYpQUEEdqREf8yt3XEnR+ix1mX3EBF
juU0yG2zAH9rnjO6jVF9HzouMS6wHa+4uMy5rqt6wvaNqPASy0wm4YQMnSRx+MFNcVE4yp3pyYYl
uxXEKivWOXSeH8VyTv/q7YIv5ksIrzUI1L/c1LjiuKGrU4Z9izp9cWUT2pnfQCqerur//1f2/oFJ
byApZ8p1ZOG2AOFlP94DWQsPZ8/ch57jqtRJhLYy43vS1aqu3U6xPgPD2GgFsI+nnHKiOhN9uVag
W0u31CVISvRQ5BUXqlNPXj1V6CtCExnHHDz9sw4TCL8b9qP+RlwQvedrtpEONAzHdodGn36TEn+H
LGPIC/6WxUGGVAPzgDKWeYeMFlEkBdbmkiz/zGZR5ehAYXlyUGJ7eQI7GlGpugnj0YoCVTbQg3Ao
8mUvWkBuyDhykB9Met35k0zsnHiw/GyvQ19sDeydXvc9tg3A/4IKSxt8q1oAH0hVQMDiYYDpEKPD
V5wL2hvv4XBumi2HO5XuOenYJuQMgnVe06X5sNVl9I0YvjgVW5HLliaLLdUnavXLesS1J+zTYCSs
Z2adJS8+UkGS9EGhtOCJAjNM207JlCoe0X5hsC6EMS/dva3mj4owIbA5QZQe2gnGnW+16mCRk8y2
9W3zg9jTNTFlhga6DSblzRnp+yvc0gK7XcEUT1ckotZOlBuPXy+Wtl0LS47j+6LyqyAPTgXeL8Dp
bCtvgO/+eeL6YPP9nlsBdfiKeTpzHgB+UkpJxk5QPN57gkQrSkwKbSQgIBR5fMFUvn+bBB3pfLMI
T56iuEKnoNkpKZtdCcANoQbYBmdPEiu+aXPgtrbFO83nggwayTZTfuN2+ULv6X5GIiPS/8/TZpTw
0dlZWIx8f37rfScwMZDUnYXpKjaIzKPjmyoAfug1hpMoMsIDUs5PrJQBY1a19FLj88ijTgnt4YXd
0AUW6mbgCStsFuNbRAqF3mcltHOC15saYsXUIBa7njJS8n1UgX33CR8Zv802jpLIwMBVUhV+KTU1
r+MHgT9mbgvfE40alqAQv5Q2QKJ3CQEQdxUvr9aL2hwT4++/qceTLiLQ6v5t+9kg3d7vfpnlGNpO
wP+QqMZi9jpDd7YObHDp+mfezi9ittE4ya46GrSvnkVbTe/IJyuPvPl2Spuc3dpJP1+ywKWY1B6y
e/BA7srlaLgUqIlrupcHpEGt1CUjWqQlPSVfM6AD8X0ZsxuD1KALVw247+nT2c4MXOXuSX4oaLaj
rPlVp4LbK9layof9txXdAZgMyUHhzPF1feIDZzA/4e0Gc3Zmg6dLjsjC2W7/dBvr5y9pOnyT04t6
5kG19UuntPVdwU4oEV9BxURjj2pq5oU/8plEay6HAE2Llv6GgXrN5Ba22DEuoBI9SeJ7aYGzzeL9
i3c5Thkc/5EslW+lV+fyhld7BK0L+9cXHSOj/a00kxqVx7F2+XIijOJ6fIkB446vxQ1tFp8OuKis
7VQ8k/xjZC/zL1kQ6p+OQYUet8we4jtJDXBY/XR2XsM3ksbu8W0VLhUfw7d9ErNddsr753rhmJqR
MZZ1ReIFRk74FPg0HzS6yI1oei8pcYS9GBnf5p6034hLOIhnfibRWbo9pO5cgAU5NVUJ4zlEwmad
mHuOkt90UFXyu0Uads3tWecEllvVn6WYrzz69EvzUOgcdtP18uQoEKJoOZOgHtxrlbFNZhzvNuIz
g7uU/jQ1pDpBPoVG9lIkMbXTyluOpZvAJuixMFwr1bLlc/dC/XwO3ffKGvtqp0Fsh0TXW6LN80uj
51DBzbhVtXAYTIXRGzWRgnXbgvyY3+46JD1xqomYJxfQgkzptAP6WanFsftuNwR96ICYKiw5ZMpi
9m0nrjs+LnhhA8PlHgR9dHBY/4ajO7v+0Zv/LtDLiwBV8dWs367qCz6MkKbjDvwqq9xQzbKMn0bG
Y/bZUGYMYMg7OXxoxoJUdBt5m6nhnSzj4xdHmj/5S+dvKi/eUg0p3MLFbONrPcNuSWB2e1UTgFiY
VcsLyJneOJZQSS6ucsxG/MzaytNwhAHiOeF4cZs0Yn0eEXo/N8NHGb+st2/TOjDb0H9crzUj3n/4
jP8mUMuWitmtD5vkCp3CVpnHzII9Lz78tLnPIl7xmdc9yiwz6GoxnKYUmwRJkH00e0nG2sghZ0Jw
9i4PZmMpXH1r9I4dD5a66yLKHjMZv1esX+7b9AEZpHX+fds0IJG7uIxt0X7RIbZQVBXG27vEwimT
uSW/3E4ljLooc7UmUc8zQ0eDfeAla4qvP41E6RXEJApWT5q/6Ih2+hFKml5eFYoC9uMhAijNn2pB
xZcyKDTLFm5aah4Jh0p5Mqixwvc24eN/5fqQRsW3JvbUiyVvxW3tYIXTE8+f2zHqIYhI9dTk7Hnu
1TTDZXJ5x0M5rNOf3YDsLcmNPH3FMr5paNxZD16i8ggDaa+ZbehAYy/dsLic1t6Sy6ErmalX6bZc
yajRNij66ge0KJagDrzqtar+LgRlzrTH/AA9EnOs2eyjuzP/vbQXTwjv/62gx3nNvzz25zF1MgND
RXkGdVCQPYzgLbnU1CP4PZ22ueImvO4za0N1bC1YMI3na3oZ2luPbEF0XKnQKilaosEcRGvRuHAV
9a1bm0xcogs8mipuRdcJfiL8gxl9mP/Nv+rZWzBuo/nTqxq8lD7A06A1bY8MiMG98On+K0g1vzPr
/JLs2WP//+Atv1WEdiDboX46hzY9w+nJKIjTCdwtOixIE4jvg2T8jslzeJW+l+QKX26i1R4w1SIF
X9j+/ic58dBoFmI8EuIgvPIc7xiQXDE7GGeKRYxqr1EfH1ex4b08LfyjGZjR6u1VsRiG0njmx33M
zThABKB/92morKVP12uQHIb1oIsexvzPeKOYW/1xhpwPdR3/PqeZK+6Yo2cG0sP7fYCIbdLv77bO
S/Lo7LJL5Gz5CR5ZEc4L9LkDrT+swGfs9MMpz1SyxZiif+3oum5jWIRZQPV+8odzBDa4p3pEd2xD
xDfUe/0i0lYGcybP2xCNICorhTeN1c/6tOsjPKrgbkrscevFPwE8EUfWAl00Pt7KiTZu+zShDkdd
2oz2zIUEEZy/4awQUoqA34kGzOXR5iYuzt32EMlF0JJtxhHLFCLc0bcJhgfCwoOBeLdEU4U6vpdL
f2bibSFPpbsRPoztyZcGsluJR0bzwImMruHzUiU4lU1Tv0cuNav009jiWEa0YhV/hgt9ZNVeNYVO
dk9Sd/lLUEkVrjlhLDI8A4tLI19tt49w9nfJ0fBvFwUm6C6AXX3B1ZNGl5lTyUH4IYeL8K48VOQG
fiKUykk6ofqEpDfvgMAz03/VqQjw23Gm6Y41RtB3icOAx/DYbzcpeCwYHfNu8ywofj7tzc4TkY48
S7NgxUv9EO6CrxlDYJWuL3/R4ERIY2XUoqqnkDUs2jfTJbFVviBGu2AoqW+QFDVBfHW+TO5zlko8
KEN6X2vFxwkcYnnUuDRhrX9MAfeoQ/MdcV+fUwTUZ52jRKH2eZpR95IsQzUR0awvHzt19IjW+Yw2
ZdWbPpihSd+6Bl+3QJjvj+zTeAOhqJkk/RlJ4f7OyfEFkKEW3wF3U5ONYGzmeFSnkKn7d+7MD4wf
djOWXoDdsEv82QZIYpeo5QGhUP+jK56YBjjGPKhSeZ1gWP7ite3SZ0T05z7AnrYHjK3kQrhjNU1w
GK/n9ZygF1FRvm+T8QVcpQHXFCJfnT+abp7PCEWeEE8TvEbgUJpJdnGOVfnWejyjf42ACaNNGUC6
VHf70RvaBt3GkNWbSUyA1nHswEoshJDRS2N5is25/p/r67+GUjnet5dG5908EeBCOsW+HxnFhotm
PpqKkRDN493vKR2rnDifU1rCvvWg444rG3XDvS/nS0VG6cvJhrJKyKuvqsMsIwMPeL6t5rRGgCJb
EfNWM2FfboNWtlpdSe47KcQbD5bM+uy5d/5O+vVDeovs9U7Y1B2iWUGLBGrd4pkgfpVBvueSnVpF
/sRq/Ldj+uOKvX8yG+N2tF3B8nBU4HeK+DihNY1rDUZytaB60hyYjAHqYXB1h+VVZf06DbLdcylm
YMWKpomfidHXUJrQ31IxFb2i0BE7rIVW0mRzwmDWKwl1T6raYO47nIKkseE6q4NzWfUezOor/vSe
JCMu7sim/P2ML8AHGR0bG4yNe6PhosnsHX6hK/9fB658z/K9qpogFqNeW3+hJGkcvVzqHEUy9CmM
52VxHOs45EmmmEx0+xdAffCRpQ5l225AUQKOi1xiXhX3bZr4yEHK+CgB0pXd1Yy+20N6RLuvhqxi
g59SZef3FEbKQVjiyuLGyWE2+OcuXyyvbObMpjgLYmMok0PyteAFXiZ95mCCINd7CvLESj13BI/T
0N2tR7rhy1Kkig84a+TMjwOF6Kig6ujTCu4j5TErXL5Z/AWAVnHTwS3VvwoF64oJoSL8ybdUJMdi
PLovRvDtwL6qPCrb+7VtC/ZjITCG8ndCtOyBx5TVXnygomQtj2RNH0Z8XyLssOOi5SUYFPQ6/5v3
rKjPyLY6ufmwfjRKDPWgelryzlYZnucPK0j7Rhm2BIRgNbugMygG/kyLgK6G82mNCDy5QpVWUgy1
hPwK6bVLdPQM0Fe0fu92gNVe828whSVAZy/13jvhQvN+00Ryg2aQqNxVX+U848yEv8JL3QAcMZeK
t7UqFDrqVpDmay6QtzgHBCZD5Xc4wS5Rz2mr7aytPb2TeLZiMcCQ3zdlre3mRSysXUZ12g6/iS1Z
ug2viql9B9mvL4M7foBqoNonga+fcwpO3tzawWuLNTpL45gvmIYPLM+ZJAqhBw7V83W8ZAUsc9ML
IXR/M89lsC50dCfBxcrmvF+S8JyVFtXO6NHOT/BN9PI4Mgk2yfKNcOi4doBcQCCWqeFlyrH/5MlR
o9TdK0I/RSK6nWaug5O7RpvlbVbTWct0ik4X76JUYJW5QgcdCDDudCG5SRj65nB3evBzXHy4fDfc
cJDbF+0NoYywreuSGu/XHpQbZh1OgrgToqiL7s/PYYIHDpKsvEO8/RE2B9nR1C24l3OWVwpu7NIi
ycxEj544qkiBZa04NDq51TAEgl22lyga/QJBNQJbTX1i+qbYFcP5Q6Wpjv4iXMmZIpwQ6F1TNGrJ
/BQXtMKPMMVAORpaiuIXs0+3FuPth8gK1le1R44aiVNKrs/4WLzUIOM5T+DJJ8mY8FdlTpysqNEz
2JpmkDRM8FvXuWPWIm4v4g6Iln8ubP2lqn44vKi5GdzXrj55Lxn3/oELeoyoOi6q2abZ1Xeqt/rO
jJ8giAwwLyxH7+zDrfkQv/z2lzDYZtitANSEhAHdpZ8yDmNW9B6BCJhEBvv9BU3DEzYTESm81/cQ
HGwWRXOCjdnKn0unzczMDaNzy8NPfUbtmS3K8mUMQZFll65s3RYYOjOCt/Svp6NWMuFlnoZnp4qc
JDiqcWgiT69HMfHWvx1VzuwwtquygBpqAIQdZ+ZKS77JipGEZWAV6RR3OuOYftxLYoKjwYpHPjjK
uNS7P6maEHxGP1EZ/EjCoffYkgceUXgBZuz/56BXCqziWQhkEE0FSmKT8nHcoPEZkuFPEeoBGxLY
6YRRuyAyDKmgsgQnG5UZdtK3cSSrQhJNZBNpyaNo7N2LOnysCWq+ggrVgaML5nI/NTejpsVdxZzg
LQYJ+DfIsigbkItl/E03wYGUXl57N7wzM75F6UloL9fQ4f6auTwITAlVJQe9h5xhwEtfYIevF0nG
WC/1E5MOQho6FzYrGeCpuCxuu+ZpgRNM0+gNL7CHsbaRX+8j9pAJV1ajtD3ldeVJvD/dBX3HUQcy
6Jp1XS1+Tu5VQd3blPwnLHOP8w+Cv6Q3B0ePrmxJR+uSjHAfM0b/l1jSH8Iikhw/cRYMBXsSt9e0
YgYkQMeKWQF8TzSE6hVGli6gtInyHWjSn3pT1P/G7uF06F9YMm01R1OseLojm+F+/YDjfcV63+kR
ihj+vo5o2hsOQirUkqXOZa4WqL7AOIw+C6AN5XywFo/8kih5JyH4USrBPJRc8dHU8V237IXAtlFa
5qMPfGplv8tCqHNgEt6uO6i5bs+OjWdgizbBkl8ohGr/y14DZ9LkDVsjAIQgJGGbqicGZXqKWBZf
SlQUNoTm6A1uL9M/SD9/KZC5KyXwESgLrB1NNNk8RRntL2AgEy3Zo7dDHyJMv1h6UQSHwnSlAk2K
te/YZh3rV661XWrHN4vr2iBobZ1+1QLDdrbcJPT9bINvynjrarZlmFhgkDoY2JoTyUfy5ia/g9WR
rzDOmdd6men/ZCOqxr7Rj3AyuKqKWBsJEt30k65qYJbwYhgJh8uqEZFJbTxLCCAU9kTRK0rP7TYH
8nC2yYpPWm9QLUduW/XY9nsh/XsBq5wzWnHAkedqyJMsPgg8S0JkioE0febgEqaUErV3OK4qZY9P
PI98tnfpN/PLMwb604DTOHxC2G0lfdLwlUcDnkumC5Fi5wN9a8XRFme//3s7wpo/1puMkAaKgUTV
1cT247QIwWk81lc/nE0iCXl+JPk2q1YpeBCCW6DOBHOzgsj7tqSmPAveYgZpbCiiUqfiXQ2r++h+
gFuxJnjyLh8A6zMHdIMuZ7lGO2sJzZ0J0RWx4zrnGX/DICsfZpx49z3b0piGjdOPzj7hACmZm1NF
9kJAaXH6y5EQNv+2tymRrXQ1IYD9F5XgOmbVDOSjZnECe0a4NAZcaDiUOMQhQGSZg6ZFPhvZb6En
FZV5kqoAUSZu3M5fp0lWxQQbfEnGhCC9POhjDfxXMm5DzOEW/uMCnZfhQ8DLL+tWF+bZFRzrGYWc
0b+v8JMDHpIXLP13V9WRD6X4wk9bioZsDI4OKBzbo1MkVLTJZh3FkzNQpqOHS+4umC5kXQIGzwGc
Xl+CPeceoXyTVNEtCDTzJVd0m5vkaPqyyx1koEPgmKXoXvVWqfgMWW1ahcHuiAwkj3tHcqApJn/b
BEtWEMgUkNuJi+FPrWd/1GhpT8ZTXjI4vgeiETxlb12/W77e0h8cJc74yMONtGVf05CbjuogBVML
Gom+Gv0P9APc6Vq+ghSdb6XIV3mv5sFru+rwNY0cFsK9WCA92IWmuD3C60OCKeAgGoCH72So6qSE
ERVjiraZWP4dr6+n3Y0ucd4PYy1cMrWabpRcJmA9EEdhP7BDjL/xHa3VjPrtlZz43QiSOiW2NTj5
tZccwRS9WE2Ffg3K3U76GjoNS+6GJNuFjiAkuDs8zGpITpkCwfWRT7aElTvNg1iXCgo11aB0OG2Q
+yJBASiwx/6zeRE7WNMPQpIE7NLgrzRH7EcFbcCFaC+FhjD6e5kL9n0tJsH2vPUWPxzgCJFDezja
D4BMCyC6Gm7Dx3HSAQKOeSV7GE8mDzB1ej+1mVb2ctU7oli+/jqfoDCNCYJX6WOJ11lS8Bx48XBL
ttpFEhVZ5he8UlQSPXdLaJ/I76LIrYDzx8fCDiOjw7gRbitVgDWzRINgldwsdJvoA4AET96NMOCM
Egodv2FMUprul9m2JBMZpeVZvcClRW1WxYDl8Pz2jMcQ3HClHpqHnu4sgha7VQfYd6OuWBpP4l6q
Edhjd+0nqGrNy5V3niu0qq91+34oAjUT+bjWZzJFijYcjiqR/jq0HLWWMHyGcQh6JRsT/JcTgXSC
aRhWIAV3N8fK7a5oMIgJBM/HpB79MWSoca1i1teBi/z+kQVKS7UreD89NBDcjxFgBEEbyQd0DHPp
zuVJnJtoCWJt8ZhLF21WnbBaeZG2zjm6XiOrMvXIPq5PNutY39YEkyMXu6zzeE+yxpLy0QIvGWcG
F3vJEcohKK9Jm6Cn953EmRg5EEfEpLCfaHw7n8x76S51CHtlJGWWYScCPKQ2v7PkeftmEkdkbIom
CJyktcLMXSH2TNV61qKKLNyq/zjoYBhZ33VEOY75p6fH4s71rlBqfOq1JQ9rGTcRjPSaF1+TvEs+
7xEJ3pU1XBGIMRyk6cTqzgvnm/QfrGGDMDjIb/+9fo/fmxOTphzlV2+EuyhTSscuBA6F5OCy9c9a
IQuS19D4mo62FuAopL97ROB7j5xtJDRQ/FrZkNRyDjXRfMmqNd4q3m6PGMaTSWftNosnlohOyQrm
hlBt22c5E1X1zbSG+GkLZ9hMCyFMdRIc17qM7iL741Vdw3ExWGJLlNpGReDGVzT3/tDMBtZsujLn
E0tiuuT55KDYJ1tdJnSneC/SxKLkGBu98eMRJ1tDCLdPM3yeqnlLVzuewhAGN6UNulwkNFRy8i/1
n0Cc+wN1ObkSb5omazSno8zeN9J+q5+JTWPX4P7h0el4hTdVd67zPPQMSTVW8dwe7v7ZAEGRvTJW
lYygRvJNvF/SyTA+HgU1mgTUZ2OYLMa3KQgqBN4b89QqzMlboLspLxN186Smh1YofiHg5GGyITgP
Z8C8Ib6NHC/Dchga6idjexpg7w7rz4lqK/KIu0qcudbT6Anl+B+iJKOG8CMk341uqjQpEAGGFEdQ
DT7/xP76wlJ0MKSW55UcofMAPV/Hh7Pqvgd7M61aaMsyoodJQKhhzeoDKs6F1d3jcrE/hz0OSHud
3whcUC7AB6/+XXp90rjYKSyIuU8M2oZNvYaiEW5oLobv75XSX7GpoAokuuprAMHHSruFOHf8CxVW
4fWrOOCc5KE/hOLizLi/etNX5NIox24eC4DWYpOdu9yvbVM1o8L/BnDGZzjRxpnd2v2btygw4n/7
agbRwk6+pDImLANoxtJn1K24crxQ0wQ9XaINhi37P+w4WZjlg+hr8GZ7b+d1yBaLou0qVWc994/N
vY6ykL5Ki/j6OKKCmBUXYlU7YejjqipwXWnuvjz3eRaQyzcTbn9HAsgmqfMoRf9zKYklzlDha28V
evlQXSyqUIQ670IT8zkNm2Dge5s5CuP+30iwwMbJi78aDO4Ie7+dmiXJaimA9ZkxqPM9RICIv3lv
e8SRR8CxOBdbA4v1ZFz0UcL5cZ/rcEXVwHJKcnPmyKN3jPUlnxw0iskVuqJEF9qpaUOCjWhTgDhc
eJ20a3V7BKCBz6uAJGtOuq6nTHE69MtXKKYxXy6zjgFN/nlYxfiJ6EJU0f8TKVQPJeqMPw7nIWZx
RZkA1krMKLjaMXOL5d0VDeLWOP2Skv1FM9oKc7aaf77oI4xdhY7aWBgY7r5q79PwaPEcsWYIapoz
oJkWAF8de55RbseQxj9WiPAAA0dbbDnnT6Vb9rC12FUk1nvTZq68z/LBgiUJ7B2Z5/p/rxX4VWV3
9HyB+nMbMznxRZNrA37vvF7PnO1rAOfUbCIbjo8Al5B8q+NHKS1qyldG8E9/aWTflmPCHCfxX/Ju
6gurs3T+ZnE7o2cS+HzPMJ7k5YHwHk76uU1+Kag4mQ9+vROhBvaSC5pbJwZzQrwJ1vptykZ6jieq
F6+f9oIF2OsflTU0505eLJl/D3609ObyQIfv8wYosDrAa9qjaMEQjvHgpIDFALaKoRWGfSX2JjIX
SOx08l9sQCv7wvEWAJ7miayUdoYIVEsUjsY52X7+n4l7BXq2Y6X5TfdhM8qFE+4PykXmOn3owYdo
5uaRf2gwPEig5CUFX8NXq3NwsoTAXZjPZ9FFd+eL18ohhazyomaY/dFme0ZMvLafk+3acQLHCw57
/Ei6YBS3xC65bGdLhEERFsCC9QAwOE5YGyI8KzNE2NlTvbtej98DqDJumRodagM7Rc76IqDzsku1
wKCgIvBAXQzSnAuvYDjs9U+bwOm0RI3b8YjatMPLh2eiqBTwZoNtbmpLdVoKRPqu6BrtfVH2Ckyq
IohN2QmqzKjRe8CEy/3G2xaCf2R2ALC9sWMZYTcf62wc/VCN5XoXjYFIspiC8obvG/tMS8+LXjWY
vOog6q3skRL8Rm63i1duoZc64r0R67av6OrNHrSXdz8G/2LDpYg6d6Q4rLhTOEUcxQzItmBC5axe
yDCyAIzRP3hdHje3nyY/0KpnN3Tdw+6N19G8s0CW/mrUtxbyvchJM2PM/hIDMD3JsGEM7hlwVB7E
oaEsQ9Prx8lfaG+S3ra+JRk2SgZds2XrZDn/dhWLhvL9M5zvDo0TM5FxvI6huSwDjcX/VQT88XdO
H8mtyo5AjkXjIZDj3oYAXeflkBXIsyNZqWDqhwgz9CN2W6EpyE0KPzutf0UDT20lst/Y5MVTlXZi
FkJJUXxmvvk9dbu6NXn4WMiLyQ2g7P0YY8npTHU4VVfULdNC6jpnW8QTbq10q9Ne2b1OuQ0jH3pJ
T8IZ4o/Ocf1E9s8+E0ofrWMamSx99QeIgjKyFZn+V+j8sP68mzwelUMxl2bOucCrfK3XN7sgQADD
mT2gvAJ3U0onnRwe2nz/3NpV7UcfTv/nEG18WD3P035ZfTVgZcMy074wJcyjy0Tdsg+aAcY8LrQt
79n+HBUwY91Vixi1jISWTJLTHVqrmhpdmcKS/EpX9rBOlqGLEclR5nvmfqxdBEs6BgLMwLoqzaeG
IpzAhoFfiWoKm25extMVFiAmsC8g40pdaWxgxsagh9is2NihrYMJhod1IEVNOjiFZwprBp/gZTPD
MAh+gVZbgW4V7+1ODN6SU1qutoZGC8xdi9f4FFCuEgxpBVM2qf1Rrfak8UnJioP8dQo0u+o/Qs4T
8bdjqWv6HpLlDNjtIOUJ4zSIwUJzvDCCiodDNJ5/PoLSpnocoBK4tBSFJduWU62TGbo95FuqnxTR
3iXcOp+GdSqHe6Yhf651oyPgfgZkI5VpkyJNZIHO/ASD1IwgmkXhcKyVwqg9zPMC60wKdC2kZ6Te
xIyHjUaM09Oh6LCY+y2wrTQ4xwsp0aq110LNYQPa4HaPUqqF4dayRLd+V9bEczNiFt1tECZfLjYo
OTiu9ASawlxZsCroZY0N6490MHSxazuGTNkp+yIp7kIhBVS38GCODncpGUGb1ZFj/RQAerIn/xXu
kTraarWbDyEKGbSzo2w9t08mYmQ1LBXxhh8CQN/hIeb2Dz+mcWeF1/4uhH/nHiHZAhAa9J02L6qn
qb4BQYhOXfYJ/mUx87r/GyTrfmaPogyV5djaylRMFlgn7EGDJ8Sw+rnKI9SM9lnWpJ36t+L2hmpE
uC5OL18VmPPUql0+haUNKRMzg9pwi0tvY4Kku/3GeUO+BsHQ/85jC1WjdpqImj+V4CoYcQ==
`protect end_protected
